XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��YsɪV�
� r�£A�\��@�4]&�r��I����l��T۱��,����$>nG���<�w��L|�����9lYж���0֡�Ť[E�Wj���K�xW�Wt#e����@��Gx����I���&~�5��U#�l�UGcs��B�k?��oN��Y���X.�B�m-�f���#
-�vƿ˩C���?I�SEl��<�M�m�ķؙ�o���M��V������`Z_��� u#*P4���P��7� �BNԆ���__����3��ܵ2��!�;9�:*
%]R�p��@�3��"X,�	�i�����sfzD��4�-Ahg,p��85Jl�"_�3#�̱��"IMR僿Ԉ�qq��n������c5=8W���������e�gA��
8U���W���f�TG�}�.;�ZK� iJ~�R����5o����v�5��f �!9������{Sj�I0|��R�6��U���^;$�=/�h^M$��S%;�=�u�O�S���)M���Р�
;�"������L?�f[��s�Y��fI<\���>2�1��ב0h��}�&�/��>�B��b���`�ɀT��A@�W�X���X��4���nXTS�Ҷ�#؋�q3��o�)1��m�i�~@W�K��.�t��LǗ�����o�x��NQ�2��l�����H׸�ƶ�nVPO.�"�]���0��ysZD���z8JrۦA��:6|*XlxVHYEB     f6d     6f0��[��K.�8�or����W�g�G�P��Ҷ�?�{d�EٔV��8#4%��'	Z��X���K��P�7E\��G;J��^�҈$�L�7O�����U2|�#D�)~\�,�Ǎ28/y'�N|ɔ��֌ׇ^0ZS�l����5!G����N��R=�}j���_�p;��� �gC�$3Umac+�;�sИ'�)Pє�s���B��
q�W75�EL�� �����P[J�$��%ҿV�>^:W����ԽK��B�v]3��Sv��c��[�e�WHs��*��[�qֹA�u�?��b�����\�J@gE�����3{�����K�{��շ�� GI94�fD>��%ƋJ�3+�����{�
���i�<m���d��7��ʼ�qX'z���L@_
����C��	z��K�Q=@����]>p	)0�^�wzy?�;�W�����7��7����u�dR��KS�"8�F�<w-��&�AʬD�O��Ơ��	��TcoIxVoR��41�μ�g�`�������Y���^��;R��b�&�g�͌�$�9_U��8�B5b3��2����/mM]��,�L������-n�%�6ON��[��"=t�xM�Y
���R�:�:��Y A�D('�5t��P��7X�D��Th������M�F��J���bW�t�[Φ6^�	%�mi��f�T�?�i�z�N���#"���E��lI>�e0խ���7>#K���H����Pڗ�"��F�@�L2�m���tlď�,�}ί�]��T�bĹ]S�CN��R�y�%��Kӕ���#ͭ�d��hX��2�U��ϰ���# �+I��������+u#�t��
m����#t*-N�+1^J��]����8���{tk%�>ςO`����}�23S�dILZ�i̖`����4yhR�"Z��Ě.=�F�=�b�y=P�����.,*I���?��nũF�ۼ���N�,7h6޼
����r#�k���B4� �#O�x?��PA*'>ǨъC�U��+�J:���;���pbj,M���W(=�K�9UI<���(�>��n|8���gr�?��D��ʟy����Sꌹt���$7�ks���'
Iu��xj�Rc32B0X+e�p	yx�5��8�ם�U�Rb����
DFir�N�|��p�2K4~iR��k����Cg�{h�(R4y� ʱ�Ѵ�8�Z��b�f�K�#�/E�2@+?G������6�?��%:K,��k�[�3YXCT����k�i�����"吕�`S�I*���s����be�����(��b7��㺢D�ŊΎqᨿЏ,ZW��iG׆��B1�[
ZY6�Y���V[�][�͌��B&�������9��*T�fuD�I�?|`�<2n��^�`��¼f �����&�C靖8N���W9 ������_zXw��j�G�.z2��{��z,���XAw9��6�\J�c�]~�X��_���b�"�G�veof�E�a),V�����֩ݝ��*=��v�\뻃������P�܎�Z ��5m��򣖿V�obe�W�a`#�f�v�sD�[������/6䨦�����j�~�L�<��ds�ӵ5*�q�&$�?�ٲ gx��h�'4m�]3#�&VJ�c3L�4���Z��N�R�7vå�򖞐�{�ì�oz%�YO}בJz�[�<ZM�2�dN��l��I�^�-@����N�]���)��%���Oc֡����֓�D����`��Y��%<��