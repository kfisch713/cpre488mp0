XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����k�B'�s��9��J7��Us`�6_�Tg��'��v5��+�������*�����a�=��-bf������(�0�}G�5����#r2還�1�*~%[��%�H8��/Gl�|�R&w)�������|i<�K�_:}�&�D%�4F^u�O�y�:�P|TRډT޼����Bx�oȐa:h� y�.�ü~,&B C���-��t%�����&�ݤ�Ck�^�$�G�uY�~�_�XNR�)����T���$�pկ��{�ϵ�����|���t,M�����c�x}E�/!�ݯ��JN��o��̪��`u�����M_�q[ks��Ƀ�i�^�pd7��[U�X�L1a�E��!�obYNm*��o�^$��XQ�D6��ד|@C�+4qRC�E�?���w�������i%%�Do���s�4�;^b�Bc�[�`VN�ߟ%$t_�_n�������߲0��Շ����8NB�7?> ~�����+_���� ��Fk�E��W�\V٥5;���q�H���V?���tGL����0�5[
�F�J��5�>�y��'&����kv�>nNr�v#9N[�/����oWgS�+�JA�H ��QY#w��</��1�0"��J������O��)�,��Ԕ��1&��a�T����Ĩ���4���b�T�"*4cD8�Veu Ґ�?u�3 f�y|��C�$���n���I�`Ϧl�+�I������.6(�_��+gO����/L��XlxVHYEB    6014    1840<�=y@�&7��]ѯ�l���EN��|�e�J؏ +�Tz����FSL	K����!%����� ��[;0B�lKo�Ih��⏳�-����v:r/ڞﳸ�n�.H��T�om2�#C@E1�ڌOdtN)}=ۉ����Y�@�h$�|wxefU� :�-z�3x�T�H~r'��P�ډ�LUsF�<?��F��X&։e���m�y�����Z��ȫ��=k�`��\��x����Ĵ_�Gd�.���	��ڥ�|�N3%���$75g�~�l�J���2��-^�.ehl�k�0&�}������!+Wq<����8�Q���4��xCė�tY��1�0}��B�2�l�s�`M�cB>|�ߍ�� Y����ǈ��������	�d�*��V�r�'�C?�V�P���C{���$����^����X�f����=]��rS�\:����!�9:\V�����Ir�ԉ�T-^f�.�9<�Xh§�o����ߛ���`���Ǡ�a\#0���n-6Y!�@$�7#��z���=+�=|a�ݝB ꋵ3�@���P��'U?2�-V��s7���%�rg�^v�ܻ&�uN��z��2(��ߛ�	�>�"�T]���1�'t����Q�>���ṳs�'+�o'EÎ)a��d �����4��pq��U����9���;d�l�]#����$��E�^��*��&|�P�'��z��ocȴmA\��Y���"X�N j�UkS�FQ��J�Ǯ����I���U_/��d��4E;�� 4��x���Td&�/��:�Z� E�����O�	�tͣ��xY�x:&�K�	`�/���w�A\-���\�AҪ�=�^}�@]cn+mC��c�*ϑ�f� h�>��Uw��i}��te���yg[x����"�;�(	�÷��b�v^��PM��!cDo1�I]!�����n6<���_�,|����B�Yq�4�1&���.[L��#_���s<��]��r�������֠��vo�G*?�7��� ��^?�!_jR�o����5}G4�*>~݌Ps�-��S���4���l�g3�D�����>��.�ܱ$�����~��Iv��5W��!�/��C cz�(�=:�\���œ�hk&��k�ES%�v6A��y�"P����ѭ��K{�`�P��H�'yY'#Kna#M�j3��~>�������?���(���%y��Ut�툅������|�뉔;�E�����4	���q��#4�D1y{�TV�,�MJ���fH�����o ��^G4���L��O7#<�H�O��<,�Fci|�4+�z���I3�qK�~�����re�0Wm+�k��N1zb��Z��l|���j`:Rf�ˬX-��rn�:�D��;����.�b��A��L)]�͊mno��xW���9=E,N�J���r��<���v�)n��V¿�^"'Y�?t��,
�:�����7���S�	���ծ�Lt'а���0����Z����!,� ���T��DTV�F���N��0M�ws���{��z	�_�}���QDyv
pvz����X�c���")v���Lu��k��F�#�c��[ ��w���P:�q�]��wg�
Q��E6��~�y�kg���K����H:f�ؐ��u�r�珋�s=8���l��V�+��2�X5/{ڗ�TJ0y����%W�n�7�2b�!� 	�c.�<	�c�M��������� Z���̯8*xƀj�,lqC�!�p�<f����B�����elÑh�
;6������_�?������a�^��W+��W F�4��r̻�&�T)#K�}>��=ں8ˬ�'���/�,_z��=u�/�ה�m��XU�H�5�)ؘ�=��w��W������m����+�3D���VOC�/O@��F����3��Y��H�O(�ABō&��-�Z�05}g��<6W)�9��w)�R�v����D�e�.������xDb��ιN{���JB��r�iT��
v�ݺS�W\5 ��x��^9��,�/��邙�VO������ӇA�Α�TH��G�'�뽭o����IA?��C�,[=j��G��� x���?Sd?��G�x2�}��!���:6N�C]��q�E�m���&7^�V�Ǿ�ꬺ��+z^U ���7eX�ڐ����DYب�IƱ���ⲫ��Z��e�ČAή�.� MCFq:�bucx[W��M4H8��X�p�x�#r�+Mz�Z�R,P��4Tp�^M�����H캜U\�	�5��1O	Ω�j� ��Ym���ȯ���$sWP����q����=�6�-�N�Ji�|���:���.C�p��"�f��H$���Uրܞ?ƾ>?+��+{�t���/pNI�a�WIk(���hF� h�l�O��\���H��;s3XC�3x�������I�_���9����F����V�אd�#�Y�y3�d� 9�5������/PF���&עA�.�hﴉ�$�Q��P��4ڟ�-�!�'� �m��ˬ�k8���o��=���
 �#Q���,])�Dd����}���̯`�+������-����r��w~��w���/Alf�'PycK�룂���Z���a�H��V�m��7R��o���Dc\g�qh_=�������Y�¥o2p-ڧ�'�VM�k
ن䛣�0_B��r��� ��W��𨀅���/臧��/��.�J�gV��,���\gD�#Mo�vv���L���-��H��\�MtK$� �f
��9�]��,w/�O���Ɏ�����`����7�VG������i��he��<Lc��5�Js�_w�~����8Ox��8�lH�,Y�a����R$51��|��n��(�~��ƫ� $ť�ɀ'�`�[��CQTsFr�2���]{�S��)��18;(����V�cS#rF
;�5s@v�Ƈ�jFH�3gS����>�4�!-`34����&�����zz�`�7�~��v�ZOg�e[	��X���-�6yy`���$Y�kB},��5���J44˺*9�{�nI�Q\U�]��]�#�(�QH(u�7�',%�k�ipư��֣�$���8&Y���ܢ�QD���rዤE�{iW.%M����[Ak~i,�i�N��e⡩��k����P��~II�w�2G>�Թ�#B��w�ۊ5j�Dc��Kؑ��L!���Yf�{ԧ����y(��R�>�"D�[��M)���OfW��.���}(W��[-Z,��w���Ȅ��`f^j��"�s�BS�A��������<�f�����9�b�[/@�D�F,�(�Q��"���#���Fi4�����1ș�É(_1��MS���t2�{�!�:(Z�0[����^Ub}�gʺf��@�VC4�w��w���������S��8 �P �dcE�5;�ɭ��A�.!�L��;QY!Q�=�Pp;��ʶ��,���ZL�O�CNY��M���B���L��e�����2�� �K��ϐ���DO��a��M� ~��TZM��:] �=�U-=��P:�U�+�E�@Q��}r���V�A$9��K����AjdEh6�%�n�&�M�Z,�	��R��/J�2^2����f~�EۘG� ��j��v��S��aw�|���sf�(��g����$^c:>/��cEB������^��&/f�ƌ�֟$0�V0�ot�o]'X?1�t����9�Gv"n.��b�9����*n7���݂;ʨv0�90/�����%�Uo�I�{-�n��U�ر���$�[޽3�������E�K�G�ߕ�8r�� px�����E�`n��9�M0�ۿ�;����^'q���}���G��T<8���ߕƟ4@Q�lf�Q�Q�jM6U�T��!��SO�7ї��α�ӄA��Ӥ�j3\���'���Ȼ�99��q1;wp�������t}��β�Pe�#��(�K����nR��+J���)�:c�6�<l1z���ON�u.��r��|2�ǭt&�Bl�v��k!~�z��q�Lh�;&̼��!�=�c��L����g3[���i��C�[o�YNZ�x�Ξ�I���pA�F�4�g尰�@g�h�����`���,��h�˂#��G�ނw��er��	�!`%��8���49�����h����t�̰Vb	u��A�?w�CU�FNCͲ��@�	7�s��,ɧ���0~ē���4���{p��0���kq�d�K����rZ3CMܧȧIY͔�P'���j�"֑�+1�R.�g�������&V��r�f>7z���?��h�86;��/ɔ=u�
Y�5X`�Pw�%#Rx�8�ύ�T�}4Qt�x�'�k�u��d��f�b!y�=b����Q,��������78�bm�(Or��~�]+)�D�xВn�jq��'���6�_���H�>o��ܸF>1��W�fu#FQ&��|�愬�k`j�H�J�kppl��0l��g��ج�=Ԧ��CzG����/����g?��#,#��32-iV�]��#�Y�"vFlg_v����=��Ԏ���v��L}�_Z�v���Y�S��l��mr���L�$�ZZ4��q��{�	C�.}F[�NL�D�H�zI��>��Txч�0�,Z �(���x��S���p��u�C���I��6D�%�HZ�8�|>xF�ީ���ԗ��h��pc��=[a'��_ooF����'|�]��9�3�U�F��*���ܦ]m�7�5:��C|NqY��9?�p�q��d��)��fƂ�,6xn3�pd҇>!��
����s�zf�'=�8��*�d>b	���[���m��h��?�@[���\��Z��s�_V��?nn�v0z��}=1�X�v�Y|�mp���rm%�:AD�1�D��&�+���<��!���̹�oc??��i*W�Wǉ�ZSڦ�ACv��ȿܛ�Kkh�ϕ��0C0�|@�D�!�8����$ShQ�$O}y�j�T�u�e���?їb���c(j,v�yV�aX�:�����6�����Zw}��'�k�,�)�-[/h���v�6�e�R�N�s�Hۻ�#�$}lx�D�[�^��jo�|2���Hײ��p�L�B�㌐�9�@~�E�4�֥Q��9O�-0Ռ2��zZct��<*���ny��1W��ꚧi�U	��)PFU`��+>��ud�љ=��ս��cX��ܦ=H�q �2�|��O��1bR���~�ҟ���R�arx0��.�f�Yz����\�����ב����<$R�4�%ۣ{�#���G��{�A2�IG[�Z�-�B�~V�BrU��
���Ft��-2v0:�u��-F��;�:	���$�D��<���u�HD'���^�~9�ܶ�4����Z��I�X9����T �`���"� ��vL~XI6V�)�)=4y�$�8��ȕ�ꝔM��b�<�|�ʒ��j�#�>/�$�f��r���3/��m?��#o���cD�$>,HD��잭m��W���9����֔�/ߔ�N�Y��66Q+7l,b��=>���1%�4��>��z�E,#8;lI
��k��nZ�G$/�4@�N��uT�l�iĿӑ,�4��|�����_V��ڗ�*����/�0pC�P�i�X�ݢ]I'�5HJ���������ȞRJ8����7��m0m���S%-yt�y"J��l{e��z�����u�����֠�D0�� g�^�>f���}\&tZW���"��%}���|,X}�|��^~�L2W��l���Z��b|z�
��S1G��bQ��� oIh�̪ቾl��(�iFW�,�X|�ؖ�	����v�X{ (�i�Y�3��F�1���>�S�x���y�;�Cn�X<k�ɕ9�<��\oT����e�]�I��FiT���6_�Ь���׫a��������G;4tc�#z��(Ʊ�|	]�����	��L��$2=-9r��;0�$4���n��ṭYd^R��'���oo�a�
D<[��ZG�XR�:MX�	���-�9Ɯ��m������;h��W��5֡�^