XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��e䐙w�Zջ�L�o�\n���}�PO
��G�낉w�$3K4�Ӊ>�ecK�^��GK�1Z1��<��^��c����T�n~ډu�d�]�)Z�Ғ��0d����}��L�qi��`�UR�DW
l��PqW����;bd�/�j1
g�����ޞ���)!LM>�E@�H��ph���t�Қ�o�r��1+�T�Ai�0ƚҙt"�̨�1Y#ӭ~��b�j��ɗ�����Ƽ�����f�!w��Xl"
^����BMQ�I4l`{�%��q�����Z"�M��X����6i����Rj.�*���R>|����Ek�4�y��,��B��.�~�ݖ�`&�'w��am����R�W�J��*�y���,�O�V�$Sn�e[`��P��@�<�ŋ���3�ca�G��n�e[�5�%T�{l )�S��8ϻTÚ� �ue,�p�sb���~��%��S���t,P�b�S���8��d�Iѩ����,O�蝾F�qT?�=`�#� �@�X��l=�D�.��2��N�z�[�X��,��@�ih��m)�c��]mv~,�7�eHmZ{�5��!b������̌�2^-�	_�8��K1[�6|�P��j��g��J�V�]Wd�h�b�ߚ�Ui�׮Qk���75���7/�s�ϊ))�@�7��n�`b�\7]���d@�Q�X��]��K<B��FO͡l�z�Ag�L�C�&\Qa�(=�J�yv���̗%���im��m�����2XlxVHYEB    3fdc    1160<�F�Z�_w]W�Q���PO�PH^'�M�-���[�LHv����s�+E���(�lk�|�$��/X��u�P������>u{������$��ETbG�p�S�tġ��w TcZ�lᘃ�+%C�We��J����j6�\3l����h!U��Z?s�.�܏
ə>�Z���r�ޙB*��]Iܑs׺��&�8v��z�q��9�} ���ʳ 鮌%!�Q,7%�0Ś���mS��Zz֩g�Ru�����k�u|~��.�َ;�Wj��j�����fW�����<{c0#��Ύ��'�`�&`����V��w}��Q�R�ו��g�&���a�}�Z���y�I���	�#hw�m�8*�.�_�z�S#�����?���m̙��Z��z(�|�]&ۅ^n[{I�R������|9b6�`ʕo��ZaB� bJ.�A{̳��Ȅ|]Ͷ&?�zH�+{�?�<�Ƒ��ũt� ����{R�NIFRc���X\�}�`��C���JRV���M�	���Cs���&XZ������8RzU�#C:֤�� 4ʜ@C����,���x9�ģ�:��f�����6݃�P��r�6�%��i7Ǻ.\\u(t?��K���ɔʿ�K�U�|������4���g4�n�ƺh`��lma�J{�^��5����I�}}��<v�ڈ�%)�M�8h.P�Jh��9]�nd�;Y�|�����7�� (�C#��4n6�.c��R �|@�+f,��֡�S�hnr���O?+�m��gު9<��X�˸#��3g���Q-N��nQ�J��sө�"q%�/��ۤ�6 ����T� d�60׃S����&�g2}]�ӳ��k�2B?��>[��dd�bw�����N���]-vd���g&?��|�#�E��1�N\s�>;���F�������#��U���,a�N7�Sc��l:��37���7��c���Q3f���`�\]{�-��3\��ie?n����	���M�o&��۶�V`�a�(<u
iڜ�j�5
Η���,~S(�Zۡ�����O�}�b�rk~���=ꭑ��/��� G���B��/�f�G��Ǭ�T�]S� N�z�㑙>)�E�'&剃�W��-�s���ۯ>��~q��֏��dY��� �u/Rs�r�|�o�۰�|-�ŜfϮ�����F���>\5��ұY�3%�j�rH"!��g<��r�M�������?{¡��g�$+��O�|Fs��y�m�̍Oz���� �~����Z�qγ�e��
VX!�V���I"ď�)�3ۂ.'��Y;�����C|�i��4p|gq���}��g9�}u��sc �X@7W�m<|}\q�{c�̰�����E%w��
�J!��q��:,�p��� "��-]��ʞA��>����ѐ?��Q����`l�#�x�y�F�p���!�]8����x����|�X}��rN�e}&��`�����:X�b�h���9�5EA��1ǝ�Ȫ�}�V��B5��?��de��M���Kg$l��{�i;�'���3�^��~[��@�Nk�x�!XM�j_h��7&����ǜ��=� ̵�.��)ඡ$���JF�>��/T���M$�*��Ml;���H^�ǭ������y^d��k��rP*���R����i�{�6��V<P-�qŀ@���6N%t�J��{�� ��`����Z�I1^��b=����x�#�֗�i�e'�Z��%�S���%G�`�f�RNH�7�	����P����sr���&�`��JM&��9%��xg�M3�{�$�1�ӳ�H�ptj�X�]7l�o6V�j��zM��00�*��&v��%�b�Ⱦ��i�2%��4�)PO�MU�,-˚!����Zw���Y��UX����)F���c�S�N8Xw�w91�|pT���8���.E�9I�\��/�V�#�XS\���)l	��@��!ک��*���#9���z�k�ҡ���T�pJ
���"_1/�[__��� 7@��P���*o�ٳŐ.��c�K[�1�*�R&�����9���$�A��.�Vm���pݣ�Ԏ`"!n���<�I�I���-�hk��ܫ�+U�X��rvY�GNJ�(	#	�Q!�;�P\?[>=Qj�k c赛H�,�zR:y�m.�m��R�"��2�O�b/$Tܚ��|�k��[���w��囄�ݛ?��T��92ݖ�z�7������qr
N��$��s�s�_� ղ��w����a1��Ћw�n�}�Ԗ���Ģ��������_bu��ʇ��5YiG^�*��2w��=ɨ�3��9x��k�\���54�}d~��"��b�C�6O���P��D��Sڧ��O��e_�C�H�ɟ,4-�V\L��+c��	����A΅�U'������;MLn���L\�[�ʃ���p���A�=̉�B��eN«/�g/����;y��T��W��E�����5��{*��� �X��r���<؂)�r4�]���,������K�Ў�}�{\>�ޡ���9ozț)a�]���Ì=��;�Y0"f��nNOtPdv�N-	L�w�V��
ҳ残_ 3�����3�y�<7�IEu~T�Q|(Mn��j������n���{�fV��S['x��� zxף�gtY��� ta��D1a[y'�%��-E��"o@��JU���,��Ҹ>~ w!��-\G�u�����	�H%�BQז^ m .�8Ж�.;�]��"��*v��E�� з��~A+�&���;͑��8�?V��?~b�TSa�l��l�q�S)1���Y#0���ٚ�Mm^�"s,��|��At����QQ���_}�o�n9�˅%fg^ك�K��%���!�%P�u�ǚ�*��d,�o�b7QGa�糋|=h [�l�#ekH��uLb�H�0�Ӝ���|#2&�X��h��"ʭ:�2�w	j�7�%��7�"H���lE�ړ�;�nH'\������(���C�yR�x%wA��U+�gB���6*���
�%��9_�f���< �^�e����|�)+z�����|R�U�"��Nȼ�"&Yy��F�H3��3��V_R���A$+�A~�jn�>'��I�I��S�u��^�`�|����$���\�i�z��Ѝ�=�Α����x���З`��u�Ԓ%�i�x*�� K�²rR�`3��8���WbV}}T��YI}��ۿm[q8f��[Q�B4,��;w|�r�D���N������L��d~�\g��J<4ɇ�|���,
a=�:"��
�:���%W*H�Gg���jz�[�"}uukv6u`3sI�]����$_�?�]pyI:�CS$Y��M�z>�	8�")H��&.��������E;�%Mnt�Ǯu!��o.zy;"��H��7��d���*�z�.C�e�b�*�f��e����fK��	�J��[A�.Oc"e���0��Erְ�`��-��F�.�2�GR�_x�����V�m;��],��~B�Z�8�<v߿�1r��M,o��1�M�B�5YF�@���`��i��D���Nh}zM�b-���8��}��iɯ�$�v�G���kJ;�0��7�1\�?�~�O����T��/��Z�ެ������2�#!f��B�_��/�u�xb�I���M�����_��wVY���{�Y�Q~1���R]�՛5^-z��투h\�f��U,o��1�9��#9�s{"�h�t�)�����r��KY�W�J�K�KATd�,�0/���H��3���s^��ցFCM8L�vo��v����u���>Z�s#�T ߹4g�2C�_�	a�$�32��&��,�g�f�P	���Ly��W��eRвޏ`؃N��rF��G���6솳���?{F�ZJ�F����1p��{��ɪ��I��'�R厨L/����y�7n���u�>
��V�c
�L�R�D��ƻ(��P3ƥ�7�}�<.��5E2�~.�뎹�l-p3/0~R��ϊ��\WP*�e
_��h�)�)�Ё&��ʃ0���� �����l���H��e�Sc�N����ek���`��\�χ/����4j9Ife��l���D���j��o�i���ӎ9Cha���{�H��Q�G���Ѓ��1<�2�YD��#����g��j�B����T�����q=�����IC|-<�T�Z^1h�Y1Q��/ݜ?�I��,��=�C��j��C�,�0�w��D9�RT���ǔzsW����om��g�`.�]b���)_�p\G��N��:�������I*�����-f��"��(��[aV 9?c�\Q/�:���w�'���