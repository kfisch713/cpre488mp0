XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���	exq�R<ZAc�|�K��O&V�Z-u\�c�O @�z�D0�hj�#��?u�mA!�z�HU-x@�xxw~����ۏ��|�x��x��	9B��-EBO����� �D�]�4D�0�B���)�7��Z�N�)-�"W�����J�6��5E0$�<c֗m��W_ �?N"��d���x��n!����|����p
�R��*9�RU҅�uwgo��`�W�w2<�?k�GU�N�m㑾�Ei� �aS��@��� ��XM=��g�!�f�P��P���8w���ywIr3�F
��0�T���<%@+�Q���1.K�Ӊ���{�������bHn懘�������}�-!e�R�ү9��tU���lQ����>t�����?q~H�h��>�BKrt�E��3�C��dБEś@����T!ԉ9�0�\kZ��qn׻[��m��QI�gy����ȳɪj�|^ԓ�5'��bip�1t�������dQ�,cI AAy�4��z"���K ��ʴ9ل�LWi����Հ��.�Z�
4�Z��`�gU�Sz��{���Q�I�i�7���o�k��c��3-!<��N���}�1���������w|��c�Ϻ�{M~БR��i�v&0�%+'��Y͏K[l���d4fM�wq��'�?�JB�`3��ce��f>+��i�=1��q�P�a���b߫MJ�Qc�� ��`���L6�f�+qqzޛ�T?��hs)�7u��H�+S��%i5MI�R�?_�uXlxVHYEB    3b09     f80�5��Ȗ�4���4ʥ�w����c�超R�����gV��$�|�f���/���R�|����	� �K���J�iC*X!�+,��!�"�#��`}�������n�������-o-$�
����a7�z
�S3PIqضx;�C�2	pmx�W�a��i�R�g��?G�*=\��ъ��M'�X�M�孫�P��)X���������8�g@���O f��z�#ؿ%"�l(�%��H�b��>�ef4u/��A%���w̃5fd��Y����I�@����(k1�1��{f����	�qR
/��N����pu!J���[���vM|�Zd��,@�����w��̭�)ę���3˘�\��J_�����L9`�l\g��d�m ~�4�Z�Nd󧭃��NtĐ1s��Cֶ'��,2y.��poN�H!�^�+|�3Ihf� ���|�l���*˔�f��@�Kr�ښ�!P�w���h#d�:*"��*tv@����Dx�_́.L)V�6�K5G�E>I�]\��[J(�2�@���,����c��[{��&l@ͧ]K���0�cH���R�`�~���J�w�t$��n;��b <�9��BT���c�)lЈz`e��vֶ#|��������3�r&��x^H`3�M���tx���Ά��YG�����b"��ᶙ@�泥"���$P�x��'ha��/ϱ��� �����8�5s��%�0�9��=?JB
9������<�\�(lU��d��j$´�Z}d F����\����Ut��!n]�.��Fq[	��?i�ݛ{�$@M+]����eސ��E5�QMC���kv�dC/g"jf��~�4C~�c
�)�>&]X�Zђ�ĉ�O7�ժ ��u�׭?�L�D��G唚�a_�Gy�:�v��D+C@)Z: D�ތsG���g�2��I����`.�z��@A�O��^"����UQ���4����(�MY��t��0;�jYw��=���c� .��ȣ�/� 8�Y	7@� ��]�z"������5��W�)7q�H&��Ft�`��x,Q�H�1��/J%Ѳ^��Oyl(5"�t<)f���� �\����������D
�����5����K����ړ]�j~
< ��*"��&@}$MW��F\ �u?�\�a�� r�^C����6"0�[�-~��=AE�I���z������P���;�'v��|!���T��Lȸ<o�Z�>�����6�\���Q��L�&h��>ϡ ~?-�\�*?W6B�W09h��Z�L�QN6�'_��Pn�0M�WF��C�k=:��E7������4s�7˂���߅���,L�dy+2S�;3,�n�^�ha��l�����SF��q�Vk�n7���'�rB
�w,��JhG�G�&nO�rD}AD~�I�@��-İI��
�� ۮ��ʥ}A#G��{{��Wk�x�q�o��ӈg��f4Aw�ɴ,h!�h3��"e�fK����'��8Xcq��\
 ��[ɘZ]_s������g��L�.x��W�3���>�#4:WB��[;Vn,~m~k\*��è*&��@.�/��þ�}q�`��6ɜc�5��Rj<1��˪����[�%	)#�n�����
�_tη�c��;�u�{D��}%�UB(��
C�U��F'�m6��\�8�=(%6� e�5N�Z�X��N��N>����
�,��oq�a.� i:ҙjL���+6�o}��e�!>NWC��^�P�N][[�����X9K�6ѻ�y�z|H��}���Mmhh�=�RwS ���[��G8<����MY��&��lx�%���a{�����B4G�56�|ƪq���^���Y�����iyA���T��4��A&�����������pe���Nh��jEz��L�C�LR� c��_a�Z��%+�M��>��	u��T(׽�|�((��b�F�����0�$ͺW�����C��k�(H��XY���ëd3�E�1���)���L y��k3.��HM��/�A ^X��u:���3�%Utr�+�H�r���s��:�v��8�e]�UV�&�uQ4�u����1�ޞ�:Y"�Nrfa�g��#4�Qі� �C�!-�^�6�|�Rd�!X�77E�O��J�!���?}"�.`x6L`���v?n��)�g,�I�1
w&I��3����&Y�Y��KR�G�`�5������Fv�T�@U� Y��(c?��A�W�S�KYk�H5c%4���)5l���ݣ?*��(�zT6`,�s��6ԛ����mA��������$Ε��B��E V��w|_jx��6t�z�ygW��ԉ��H��W�#���4��l5%��<c�or��^����!�Y�T(85cݬ��i�*vt��e3�\
��%Зm�m�ʭ/L͈5x[�9����:���L�*��g�]��<Pv�ĄR���j�ӥ��tIE�/�?��:�j�>�o�l@�0-�~e���ca�I����@���_���!��ݺ<7�󡭤u n\5Z(N�֋�d gp�Y�:p�>�����x~�'�?��o�"Q0׭�T��m]C��ͱ\��n�Z9�]���w>�3��T��yZ�U�Q$��hRfT`0>|�E��=�3P��=C�����;��Dbd�B��j7�C�ir����C`i�������=��h�P�/��26����k'�ϫmZ<�M�Ϡ�X����r�i���ë���mmm�s�"��gMW'�a�������ì��w�S�#�ϧ`���h^D��%1�S97޺�+�R����F�n����T��r|�����:��u�ެ:\"��
�ڸE1}`~~&�M:���r�]��F-c�M�\�ߵ/�|K�k(+�q��E\�Q��E��łf�_�$� ��F�F�~n�������5�J7���-.�O
G�O�u���ͥ�Ͼ����F���+/�,�qǥ�݊���E�@s��ht��z����{�~ˤ헃�K�Oȯ˲D0��d���4Ɍ�w�oE�A +&e4IR�1�_~���HM� �	����K�b��զ���l��� ��2e�>��W*�����R�p�K���	�����$���lp�O���ZWE���m�\���Y��K7���P�o���+Tj&��Y}�L���"<D�jk����	��>�����](��4���g�O��q�<uYV �qҤ��E���J>氅h�b⿄"�2�{!����G�C�8�mX�8�|1�C��Ú'���gp�)J��a�	,�Hp�
��4M<K7�� ���G�}S�u�?u�j����"H��@kn���"�Oۊy�^���.U���M�;gD �g�<�@ە,~�D���Z�5C�BLH�xL7�聱���	T��S_���� ����q�{�W�=Ş�,�f�<���ʔ¾�9m9t��1�Z���a��'�G���x^��'��kճ�ڳ�*ZhP���7�R�Seێ�m�}8t���k��/�@���+Lʥ��D�x����0�樧n�]>�lA����@.N\���ނ�1�w|�;"���s�L�����5�O�Fxd��ES���@�лCdy��[�+�	^T�p�F�$r�99x���i�UJ2���asU.Y���:}}*��S� ����X¡�J �r����"3�%Y1.4{1��N����E]j��͏�x���ť��p��Z��~&����q�Vhߜ(j>��H�A�j0����_�.�(0{ɋ}H�4Q���~*���uJn�L8k0]C��+�1��΋�x�����~v&�hcŊ٤9
�zXo��2P�u����c;�}Dͳy遺���-�i��D�F�F����4�W��W���nm��Zr\m�[