XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���M���q��ڑ�47'���	�Jظ���L9`�=�Q�R>Yh`�]�у���^����BC�#���v^��x���ET$ �Jx���J�Ր�#;b�p+�����/���� ���R0/�M+�lo&`[O�����w:�<���%`@�����λ8ѫjk\dg��m�K淴�����&jSl�tV�HE����G/�-$K�nIu�r]~��l��c���$吮���c_����F��Y��mVK�yK�O����8�P%ّ�9���vg��V{��E�\U�kp���x�J�΁�`��-<"�S���Lj��s�QO
��qN��f"uSՈɰ��>�&�\AF���:8������1�cP����=�v��@����E��lt���a��(놺.Y�=�%d�����O�
�r�Z[�H�J�QCq@���+no{�-%`T��(�Ɏ�7.�����Gk�yf�qɌ���.���/���|�SB6ɾt7R��3�9�;Ӷ��1�����n8�p|NOU�p��􅩿��y['��]��c�C����`P~

����L�u
��q��_6�0�_ �LU~+����n;�;��v��Hh�}<L����mtK�\�x��5+�b����H\�v���	L��Ȕ���6�즷Cй(~h��i��k����ΐ{-���h2N�uc^�LO�V�*���%ѐ�5�uu�������לF[ ~��9�V:ޗ�*�U����UQ��b��T�2�"L��GXlxVHYEB    dd8f    2160�C;�zdX�A��@@�\�M�no !4[XT"Zdn�����=��V@������$��|1%H���R.}1��w8j�>6��t���{��}$�Ĳ����N��_���4+4�dz�^1��>�Mn���ܒ�ƾ�� �=#�\{�Ԏ�]��	I�j��ü�O��W��돈g͑���}�;y��7٦A+�~P�G����_��ݻ/�q��5�yB���
0[꫎�%;0}8� �����nޗ&��/�p:4����MH���\[�{�3��I�\x˯����_�A�^�3kt�@9���@2��B����RZ�����7r����K{����l(Zƕ�L��Y�c��^�P�g���I�&��z:p���ί�`v1:�t�f�ߚQ�z���^�_��U͍����1�l��n%���@��nd|Ac����.�	�Ȍ��͓���iĈm���J�}�����4�Pz3,x�w�:O�ؕvU��x-K��2��|x�\�ѳf�����e~z\=�{����?]�+��s����U�':��f��!q��.�h/'�;�+H�\u}��!,ڬ ^8�y{h���%����c���-���:Йz0�l�o9�����u+0�6u�r�m�L���x�%�����W�0�E�ߢ c�ql���}��cDUP�ϙ�&뤕������ �\�ps�5
*��x�N�&O>��}A�.��́��Ȭz��p�A�PSw�>9�"��T*a���"�K����\zI٦ų����k�n��9�����]&3���u��sN�($g�l`�]�|�2+�"Ct����JʕP��%��,cO���}�'��΍zd�W�
	�m��	���P�{~E�~��E�W�C'�l � U@m��8������Ǐ�y�R��8J����H�s�����-7��V�A+5��2�$�?�==;��"�CS�w��z�f�PSf��1O�M�.�-]�F�u5~}����Yf@ÝS5'ԟ�eZB���W���;ztg!Ԁcz�������kk���N8�UVD�݉�$�{�f�D��9����dy��H�-.����!�
�Ԕ��P�M@�GZ���(tk����_F����ʠ���Ŗ�@��SͅM�Q־J3�"�!�PK��@���"K>���@w�"�� M�I��UG�
y݆��X�Wu���>MǺUr�OU�Q|�q��ջ��
.��5@��e'� �O���"��8NSȶ=�rD���ypR��MR)*�iǼ�HYlp[�0�>��{��70z>i���?m��{� ֵ^{�I͙B�ZgDG��˝��B���pK'Xͪ��1��A0�n���������|6�S�o'��B^]�#xZ����c{�3�h��Y�ב�h�z5�2�1_���f�0��#��a_��p2�����2��W�������A4@S3#W�(N�����"����^�k��fY-�I�������+�U��8,A������Bm�@���(��,�}%�֨�1\IK���R�t2�&����hBn���Yҹ�JO1*�gB�b�8��I�cs�Q _L����M#�_;�y8�ں�����bK�Agz���uq�4��!~5c���،�������6�~w�2j��8�Y(�HB���5�L�Q����&�֗sECP��&�_^)�%\9(�"D����*�|���A�ߎ��= &��������CM`Y�x�_�`����������Ak~�f��o��|���9�P��g%qvxI�_);����U���}�6w_�;J��"�����Y&ʹ��b>��fbx���G=^�L�� �U����2�J��cY�P����p���rV��sB�A��%��|b�����
���`K�~�ѥ�'��	2 \<�/H�?������>��C�b$s��n���t�q�� V�$�������]W6��"� u���X!��?���'B�_P9c���nO�3u	���B�=��N�*�$;�hb��{o�5^��t�ȡiN��b���Ј�(A��W*�wQ=�,��:�R~�d#@[q��U[,��VU2>Й��W�X9�]�+�n����U�s��Z&S|3u�Cۨ�ٙW��$�~�U�K�u2�ѶS���˩h�ڲL�]�9V���Z	8����sHz{ �a�_�gט�U�R����wZ���טs(`��V�o��p$��Yɒ���5���~��`m�l[��	͔�ߢp�d�,2+AR����f<�Tr�+���V��7|�ci��
�|�
�;������zʩ���g��.�뮖� ;��ԋD�����w�i��E���Iy��*�1���մ\����jz�tj�e�V|�0(C��훕�M�tƭ������v��KN�9��9Q��"���y4�2}�8k 
mm�"8ڋ�NQ�"[
O������b�M>k�V�˨~?t�t��.۬$�0�,^a��{/���A�М��a+fd�Ղ62�4W(�[�smi��S�=�N?�%D���Y�  �(S���0�;�e��$i,0`�g�.���U�����@�/^��M"#�Į/Ⱦ�`,w$�]HI ![��냳�o�eU��c�&C��p��ej�����0��������L���l���>{�1�>���md~ϱ)q=�81����`�$!����K6;��"mш���1�p�qy����ƧV�A�ޅH�_����V���h��I��������&h[������ND"���K�2��$����(z��a�i�DTJͥ�]8n��xTF��Y���V�$��7���ԉ�DO\ R�C�Ȩ�B?�L� ���&u����=z`2C�w�X&��1���M��]��_�F^�cȵ�q�M�ah ,��F4��e�+���1ٽl�qF�����x��hrx�$������=ظe�����g(����0zR&�P��s�������W�Fh��=Ǖ���g�%�ıf��3���F�70�ih��B)幺�A�'|G�[�7h�؊���x�*�!�L(����b��cJ����/�/����
>��R��[��0Dw�e�{"������fX�� �ohV����r����7\�u����4�PO넌L�:���q��ۥ	L2�� q�u6�qq��K��x!)�#�x܂b�h���(ŋ�%nUI��N	G�ξ�]Zߝ-YJ�']��p��<��I�LH%0t�Mߪ��E�G��u{�v8�ٽI'`����0��M�nd1�����b���`d�M5'���Lj�Fvƹ�1U.�Ec-����N�"�}T.�E��3�1�f������0֎���*n��
:� O���W�G���M��sjk����6��Q��'��,_F`#0��a �"w"����I���A8���=�q��j���mwB��T��������d�9"����I�9SE�q�T����H���8λ�� �<I̥�9^���z�`���?f8q6�C�o.�������"�%�)��=/T7:X�w��̛R�#i��i�T�<�+y1]�+�M&��!�n@y��ج��oX��lL:�K��ѿ��3�E��Ja�^-��QJiu+㮛��Ycj��C;��8���at�vx�z��6n��M+��01��s`�_ژӊ�ks�wgj�ċ�~L{���A9k����^2���/G�*M�F�鴕E�&�Z���x�Ap�\N��D�t�Q8��c3zX� ۶9cҫӠ@��1���@��}��I�RG� �@�w��	��2! �-T���'�ky�*�zW?,H0p���z��%�9�����	�ټC��Z�l������r��N��A��m�jH��L�Ms$t���s��n�.ɱ��~�<*�� ��yII�L�`�U鉍w190�o��GV�R�^-��\��?T��a=e�v�Z<��ĩ>�D0S4?��0h�qQz�D��ȿ��tI��0���DY��(;2��j*�2O�b��5=L����s�<�=��X��x���ҎO��w����Y��Zc�7
���yuQ{�k�H�D����ݖB�I*�_'L"�a�J�Kƍ�������A}����K�}�蟅�p�g��J��F�@���R�Y�|׊�?���1WEHZ8$�k�5������VM�5'��=��h�D\�0=�ak1�<5�T
*ځ��'8���I���ϵ���k���Yc��k~�%Xt8�nh��s9w�n��S@��3���ò��n��k�2x�F� S�'����
����he�1��,��`�����v����Y������n=x�Cy���Ư����V���J3��d��]�|K�v��J��S ϰƚZ�z8��&kě���-oL��ò?i���?E�z��4V2,�F����h9W-M�S�b�o7a ���zo�Ps�f�9�M ���5�/���pSm�h!�ﲢ#���eDQ��[a��=�?��i��/�ZΏ{�oI�͹�C�`��{��=���	e�$�>aD�n@N�nNm��+jb���6}@��2g�S�|��_f�jgB�zq�7Q3u2�Yҭ�Q)���d�91�љ�,�7�  �b%~V+)���p �����wv�W����=j�]�AiqB6����m���+f%�ӯ���*	�a.�� �+�� ����ĞHsQ\дC"��'#A[����A������b~M %�ScOoW�â�&<�6��C&��wr��v��.�ef|@���'UU>[V�Oet�H/�:�S�N|ב~lE����HI�1qzp����*܈,��6[�\M����g���(tI`�r��G�Uܭ�0ΐ`���ؿʉn��nS	�ַX�fպ>��t��E���$�Zr>�;������0��Zƣ8�`�_� �9M�����sL�[^���<� m��D���6��"��ˏf��4�>"�9�-�H^"]$�)���H��@�<qxR�,���lRL�����lEv�yX�x2��c~X��l�9�C@0а�Km����WC��6~��ڲr��֋�㆏��}EDqZ�F��{��m�x�|��$�U���q���=u�N�܍ ZdqK����:��>djSw��)�.;��#6`����
r����&���z�W6d�ݡ�u/�J�d�l�\v�8.���P�u�n9�99#�JQf�F`��=u�I���.�K��U��q� K��I�z��0�Ĭ�ps��(+�=k|�jtRI<�*�՝��IG$[�����1}�uV�9c�~=b���"nN�"c;H��<�i��|i,�&4zjGm�VV�-��IJ61ʢ@��������wzMw�3���o,�v�#�y`�b��m��0	:��|��x1���kʑ%�3���"Cn���x��p�я78,Fk���sA��f������ae�G߽ț�7풅�KjYĻU�+�"d��}(vy�<�m*�	�#�F��G������ԅ5^[�mF����[s���ۯ��@���N���<��X�Oײ
����������N�w�ۅ�ݽ~3�n� ��]H���ً�&
�&V�Ov����y��&�V��T�zE�&:a�Q��5uk��ؐ��x�I�2��V�i���\\����/����,ڧ��'y�׼6��c��*��Fɬ�����B>;yR\����Z�}fߦq#�ѳ��p�WU���ᒅ���6!�|�z���;�2fmu}ޒ�=�ާ"]����4$���}��d�\e8Ir0c,ڑ4�x�שN�Pj��Tz��ͳ��y��}
I�s��z��;���J�)z&j����p%l}2���1ࠚfح�<>!υ��uA�aC�/I�k����@��)�Y�=�W�Kv"���!@�ؠq�@�����^q~b�����ƅ�)��\���t��0����Ec^�m�n�u`L�:�0y�a܃0�"S�ښ#�կ�c*��W 6����s?x���#�9P
�<
���j �Xk���+w�^�
z50���Js�Np�=-��XC �H�4h�n�`�~�Fd<P-��e������!���>��LJ�+�C��{ ��b����|�h����!�U�`�兖^8��(s̨O6y�*�M�߆�D--��<E`5YZK`:�vuRZj!����..�q'�!X�H2������h���q)�ZKy��}��oL�҃���]bc�2<fk�g��F����٢�f:�(�P�S�}�y�
�:�A��7�
��c;P�ξ)|{01���f-h/w	~�	�͚�g��v��i��h�ZCl�ȯ=XF���Ur׌�:T'�%s�C��i�)�8tcV���W���	�A�
(Z�m����s�X&�,�?�t	=u�V��ٸ��v�q^�ŧ�?���;�G4�^��1AsX����؊�$�y�k4�}t���:#I���e����.�p�f~�����I?��ta���EH� (�f�#5$�U;�+o��@FD�u�V�),��@�^�,=�O�v�L��ng꫶M��UA��ZA�L����M��vM6f�����m�Ӻ:?� ���=�������P�
���Ap�b�l׈~c�E���%���*�
^'o<�h��ӡ�֤T��;Iw��y��J0�{��3��hfZpCē;ĺ�/עa�!O�p�pJ���@�(���߉���#�C_� q�����R���kC3O4����kX��M�x�.������cʫ*D+nGB��N��[Aښ�>�.nC�0����D�D�մ�V�����9ˤ�=Ȟ�x.ee[��LN�D��M�P��A���B�n�9�A)�9�~̳��HM$Pe�����A��Oe�}��|�k�w�6%~{+8�)�%<q<'��ނhA���!��?��H�O"9����i��&Y �J�7��W酜s�,N�SK�H�Ю~׋}\Eⷴ�:���p@:��6�m�H�����3}(o�5�x�g���8�E����:p�0����߿#��bD�LM�f��-B(p�4Wk/�i�IoH�h���KS�}�U�q�ubݙ�ꢬ��{f�C|�2`�Em�����z��kȹ���[(��8�,޷O���Jp/qP,�����˿p�a'�]�ٮ�r�H 	�ĠUL�1��^�e"�v��Ѥ<rW�	~:r�����	��G��,P�5���_�@i��
B'�+�Q��M�g��0����CG6��nd�ta�-�i�Ii��ݕ��xo|Eb"�5������Ys��Sfܤm2_�@w"�v�g�����P��s��8�\J�^��e�F��&�d���_����N�SH-���{aF�V�^�K��F��������t�V31wt�[fIhs�Ï���UlG9����L����wJ�u,X����1�;T�dZi���f�K��m��Pz�l }^�%�=9�s[�W�@�)�,C�A���*n�����st���0��H�<�d_'�8�M�@��l4ow��b��K�97���i����b�٘ءaV� V�Kϱ�	`�ѕ�5<�Rb�w�'P�WsXb�.lJ��vS���Cq���d�\�6���Nd�$f�P�û�&�0?���W�c��w��GG�2���-}g�A��L��HW���W낯!&��v�(�\��A�a�]KT����7
��;�jat�E�f.0�x�G��{���aw�Hc}��i d���k�t^"���f.��r�C҂{C7�یZ����8A��c�9&~���6�����YF�a���>�@{Ԥ�m���o�}��f_C]��^^M��rk��5Xk1��ͯc|XN����r�dH��dŐL�Oc�{һ��M�����񐍊G�l�<�d��3o���
+����$d%\3A���Oˣ��\�H^�!�����������E^l�d�
��;�)�l��-�uZX3�Պ�D�X� ��s�$}��")�!LB�������ٞ�3�(hx��;����		Hz���z�\`a�~�����K�V[��i]JTN
�H� l���J�n����9#8$�t+C��}Lʤ��H�y ګ���$��!�S��ʍ(�.����*�zקad�<�j�$d���)���Ẽ�u/��q�(�� �=~��T�����Xɋ��8D�.���0��@Q��f��4Ծ\+�N�k���@n�� ��DO��ylw�!`��g�3.jL ��(ՉR[�fj��ý�v�SZ^	syg��פC�I��m�L��V[U=ޚꃒK�lȟ�@V�f�ƵEQ�r%��w����� }5�C��8�o@`�c��$�-���@���~D VK3�u-fg? 
)�y4�r�E4�
(��$��^T]ڬ!zW���w��2�*��]��\v�����4����[k�ӧ[�#M:B�*`�ǒA