XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Q��ؾ% ���W�Tc<�*�R.�8ㄾ�cN.������[>T+C�&x��&r#mހ+M
%���F Օsys��\��
Ў�\S *�֌&��,��-v���PV��MDb�
8,Z[goX喹���GŽ�L][���qpN��d���4(U!e^�a1&, l.��o�O������a�
�g͗ZLrk�9���ee�**;����:�0N�qKyWG�
�q�=�s@)7Z��ٳ�<����� �k��9���$�_1�4Z)+L���c@��ԗ?���t�׶:�� �
8�� �;Z&��9�ʵ�-�(��D�xa'���Þ'��&�Pzm��ɚȀ��r�����i�w,�O��g�+{=�؀�;��+�-��6�����#c!��'w��j�GFdy�,�˛�Ց���3�*'+}9�ͭ6�+EK�q78�캳W���
C�˶Q$�!/�F�G7�2�ƒ��ņ��+��+B����#�/UVE�Ɩ4�����]�b^U��ypN@��Ͳ����v�Q_��|06/ԕ����G�L>���\=f�'_��[�N�P�Z�qRoo��͏�W6�
a�?����D�凑ɺ�A����3"�iOQ�J�H��5e+��]&��\�Ĝ�SF�h�0���o�}s\�RX�d���r��|��o������Q�0q��l:����5�+J�3n�n��z��";�(c$d�'�X���ˠdd��mE��`�%�;�8�:���r4����ګXlxVHYEB    3b09     f80�.�[�kܷ2�O����j��x��s�pY[p����)����u�{��]mFj?�oV�3�8�Q�^�ں������-L��	<n���2i��"m��&#��o���φbX�J|��b�k�4bʝ'��	&��Z���8Ld�!��Ez�EH���Y���A�(����l�Q�R7up���1���0>�S�N�i"p���I��ό�[����#���<ս{Y�J1YHG⁑��ǖ��k3]I�f[l���s��A�Q@��V�kÅ��9"�P��̲ť�tJ/�Rd"��}��۷�`7=셿v�X�f����o��0���1l��}_5W#�!X���?|4��+��t��K�d���G�i�u��Լ3eC\_�u�p���ꥻ}�&+�jd��wM�6��Xإ|�'S�r���)v�ύ8?YRTA٧� ��N�X�Ϋ�(�n�ӕ�f3O��	��KY�r|�i���3�zL�׿�wB�e��#,�V���;�U�,g�*B�^2d0�{q�)�C��1��.�,bl��k��T]v��GM�Ԣ��O@�H�_G3���:��&U8�h����o��@�)�$����W	�w]��V�q^����U��c�=IM:�sLFnr
=0��T|͎�>R�=#�O�����B�`*�=lS\��K��=h�:�&NE>��;}\��������e��]*��f��Y����Kce��w�������*O�g=�&p�4z��?�TBY1�ܙ�*���P�5���B�炞1�y=�e��n���۝f��hng)߭����ۈ�,ǒYP�颥����pB^(�7b��x����dB���H����p����0�������W5p�%�q���(��QO粳���^-ٺ��b��u�V����� ��/M��U�@�9��˾���0����9�\�M�p���<s��kE�����@��0�}lw��A>q���6���cQ���j20C�4�nn�A�Ap�Uc[wG��sSC*K@(�K�H���~�1��,�$("b� �+d�o\O�5Ɛ	Uu
<��(�F���h�l�y�)?AE��0�`�imn��W�W�U"���z�� ?�#TF-l�D6D���J��
��<��Z��<���T��Z��^�I6��W����3s�M�N�,,�U�G��&��l�rK��2�����K�&5�xOˮē I��xץ�G6T�\�˟�<�d�m8�:3_L�kA^f8^>;6Qr���ඉ�*"z��RijR�`�^V�`��El'�#uSYC��R�����r�� ��ou_~�����T�1��l�jB�6;�b��u}
�\E3�-�6{�x���~6h�R�5FTq�
�GZ�&��v߶�g,�ˮ򢟱 ㅮR������]�>6M���J�'tV�$,�t"
ś��m쿛���m^�A��X���y.��� jQ=�1��3+�$A��4k�B�e�-�~zK.�˗�N
7@DO{��K�DY�NB���������xFa�ə���Ι;���6�!����vC��o)�yM7rg7�'���OE��s��PDXȿSj�����r���*��"U�m�g�����o r����`�p�����G3��B�R���3-����,�w{����{,���oѝzS���,;J�ɜ��F��d��p7�@�ݪ⍪�:��P�������7�s	/w���8��S���6�\���� �?^-.�E-tҍ�ߜZ�5+on�@o+�An=LC��e�M�M�J��!�sV�. O��J`�K]IR�U�\���-v��>Z!���[�,������Du��S����c�^�������t?�Z@�У�H��o�d�HV�Ib���b�3���h�E������ۑ:��k������,V�LJ���]H@��ߊ�)�A4ב&�?4S�Hk����&q�Y���Q��4,�`�dx��,=|�AJ�^�U�,��-#�xhE��lR�w�|3�F���uk!t`���t���F6�7㿯t���	PZ�aPk0��dd�	x��>�ߏ��A�;D9Dyua�m��ʯ���"�
�C����`6��V�4x�/�K���᷺ɱ�Bq0;���6��@�ιKt���s3��*c��IQ�J�z1`���8#�w��hQL٦��ʝ���7��\����Z���rJ����z*�ua�Z8�St�6��&$G�k�J��F�,���vÔ�����
�o��o���Z�f	"�"�>���@01�3(OT��Dm_��ذ51j�<������e���\�� B�%Һa��ȵFk~ȃ4�MI�X�\ʗP_L��Dwh�xV��o��/ �r�ۈ	��&�|L�V�S��Vf�������?��6y����x���|%�ȣ޿̬��2 ��w� 1��SRH�i�;42��8*~��9?�K�k`��"��LD`�q��H�$nԼA���7���d��[�U�hI�8����ٹ�]��;���{ �[�T���SSb3��.ؗ^�8�
�� ���K�o�ct�;����~M3�;��y�%$����tW�͟�ʪ����o�D�V_3�&�� ��fn0$�U�8�Ck���IO�����C�B��e����7���*?	��!]�+k�M'~��\�xk�I�	�]W� ��R��_qk�����w����{���x��gqO�&�> T�~"��)2'�=n��%)=N�oږ�D% �G-�ׇPc��o?�L�R�g򯌿o3�A�nő7��J.��%p�Y���y�ժc���2�k)޼,���x����x�3�w!vT�n��+>9@8N���$$̾��c���'��
��а��̣.�q��z��
`�$�����W:_�~��K�W���o����;W�4����-�@ y����������̜P�� �Əa�����Z�t@8�� �����k�8�S=�� �Q�a�(���j�R�]�M���
'�!b�Ă�px���?��W�WS�v���]��0��U��D��}ѫ�{�ҵLI�8�PB��Q�j�=-�C��k �0.�\�����ڝz��W=g��^��V�mFδm�������ɰ=� x{��j��
�g����l�@FO�.�Я�}H�H����jߡ����z�i���8�a�5��<ή6��A,� B�CNN�q��h{f�6�r�����q�tб -2hs�Q��c��O�EMVI��?(B�	S!���>��V�s
�rN����nq�!!�`���N��;�0A����Q�ːv>W���Z`�D�A��6�QX�9-O�c*3��)񀭡�������C"���k�����Jl��c��Cˮ ��xk6CJ���N/f1y�AK���Pt��v*�ZD! U���?�ֱ���ɧ���w�<�Yz�� ;�ͷ�C��s��J�}�z���F[�sX�伐��"V�ެh2�pB��E4G���i��R2��]��	q4��U9ׅ	�Mgj/6)f9*�	�<���Vػ�����B]۷��n�v|[O"��oй���ڋ��r�B�����!:������ˈ.�ߏ#�P�H�9�Y�N��\�F��\�㳌V炂��[�3#S*�~쳳YTt����fe�W�ʒXuz�m�p�jArK@,)~�����5S�s�I�{tv�vanY��UkT��3�o�����,F�5�Gk�i�u@����쟙�R�D��i�D8_� ����c�������x�Z��e��b��J<]�J ���#��~����P�U����ߜq&B��0�   �2��)�c�sD�daoL��<��0&��a��]SF��@�����T��_��W]o).�'z�$*d���/s(�}P)A��&�� �T�z(ri8=Y