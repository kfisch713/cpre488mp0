XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������y�JO�p�&U��;5��U?ca8W5Q���#zC>���42)X o�!-��*�jw�ș�7�v~�00���v۫�y1�ЪQ�	�q�cƤF\���Al��H�J�%}1$����uD$e���F�����)������H�:���}°2�*�zƿ�D�n��]w���a����N;������PF�V��{G�$�	ܬ�3�`�� 	R*��_p�#�bz�<z��9�]�8��q<tS��1�%j��hb>8l.�x(V�Ŭi�|�+�s�BLm'��ؖ���o�խ�R ��>\,��O3x�UA1��
�k�������dٔ�n3H9M��8�UV��+�����O�޺m��/���r�q�F��B�w<M#���%Ѡ��S��`u�P��ZP�/�]��U+�0g:<���fp,�Ox���}�s�G1_	-�1���nNT*ru�7�-�{=�c� �&M����6C�%��f�ɳdf��,r���G��<0�a�^+��gS�c�Nh~��&k�}�$D���S���V$���˥-l����*L��Q�^��D�#�,�8˽C�X&PΕ;n�y���\,�Wr��ӛ9ʧs����q���+�
�-����~�֎���]OE$������<±rOsqrN\���~C��K�&�l��I���kp���Z�������iX�&��z6��P��g##�:�Y��2Aӱ�V��d�畷N����,0��31Ce�����4�Pm�3������XlxVHYEB    a037    1fe0"��w���愭���K�JHc��P�'�G��F����#U/X6T��s�o�S�C��1��^�:i����'��U~KA�,&,�l��.�Z�N�e�L����$X�8o�u�N�0-f���v��w�s���)����#0;��N*O�����)�Z�w^��J��J=��C�H�ϒ�����<�<������j����6!��j'���R\L��
�K���D�)�Bc����M��gl 1|���;9:x�3�. ��0M���S<�H�ڹ �ϠԴ�Lڐ��c2�{$R��b��"��^�=:3ׇ�d:6�łZX]�hs+B_$����r����H��'V���=�cuڀ� Ui$f'E�|IgW����Og�`����Ȫ��ZJZ�O�겨V�vq�����R���~s�Z-�c�%vőU��κ!����ن�� 4��5�ϔ�K�;2�cʦ&��gm��$��c��}�.�/P��Vҋ* f"q%Y'P�$�>Dn-�㬾��F7]���/7^�
���$a��"��Q֩�A���ͥơ{*�7Z��9���# S�����;!��0����� :P����[?*zf�8������09r� B}�^�7��?K�� �sK��6�l!�lL�G`��^���g�'0G݊�)V�H���I�����?�RqB�S���s�'	%i!W2���t߈��3ғپw���)���p4|��vNk��ZE��Z�e>hnc��g�����C��By6��9��G��{��&IL��a��a�l���=���Tha�/q�	�~�D>����[<�K��s׷�5��2!㋦z�nD!�5w��2�ppy����&3c4�a��Kux�Dj���ġȀ�=��W� Cͳc�w�m�=��.��0��w�W��/��}��Jȩ@�`_#�����,y��#"��c����a��#��N�B0�����ǉcaN��/i4NB�&��D��"Te��wKS�Z�z��B���	�����Pޱ�Ȫ�P���Ȼ��C�J�Ś�=~5k�`>��G��P��n0�xDk��	�	�+�����B�v���q�̦�Z��	��Ce�	מ)N��ʴ��of�_�/��'q.��@�j�:���}����_[-���QDpY�Æ�o�D#-�oD,Z��D�؊.ܗ�-7� ׵����v���1Q+
��]jͫ>!��T�XWM��\7�:?��h��9���� ��t��v
�,�E1)�������%��=�����:�ߣ��Ȗ)'����MW�M8����=�7��5�V�1\-/��� �y��#�<ا�lx_R9�r�,�~u���ϡN�/�N?����1�0��^�̧��`� k�i�3!��Q�GSv�-])�s�.uaF�C�^~��N9��{q�)�w���B�/?�D�ݘ�����D}�-���4���3P��Vj��#�H	ri�Z�0C��ˏx�j@�҅���Q\<|�����7�mc4�����#����8�CH���Nm0���e����Ԕ�����[2�\��c��U��{ֱ�K���
9��qebIr��A�]Ɉ_ �N�;�_�ޅ��&�:�']��,i^�����C��}�$��ݠ}c9Bd�xժ��]�R[J$�C$O)d�=��yL�_E]u����-\� GS����,QO�&q�P�#�Q�7:aH��'�P畆͎����'�(�vzWR�y�^�`@��;F8,M��>S��=��Qi�A\>��B�Z��t�dOE��J:m�ۊ�+�IP	@���̚�f���]I���V{�Z�睼tH��}2r\rBr>�i({py�1���?o���W�16P�b��F�rM�2��ʋ�5��M,;����[��R�G�lEy�w5��$ꃨ����8�Q�U���Y��/��8���ߌMj��Z;4^��Fͳ�b�b}�n;��m떍�;E�
�Ud1�H��Q�jpߑ�v�`I_��.3�۞Ӣͣiv�W�xw�������wu �lEFqI�x�q8�9���DMOAF�;�2C��7͕�t��_�϶6&�1!YS�[1�4%���{�m	��m�x#0�kpv��:�\�%�8<n��
0O��%ơ�0�"j�f��SNU���_ż���Y�U��ޘi��~bݙ?�����3 ��;L4��vD,Z�ix�cV����-UJ�6����2¨
���r��o_�ɚ��f_]A��{���Ej��6G`H�jx*q����se
���磰~v��fxh�M1����o���u�'�	L���3�,j�'^�Qﲈ�בpo.4MW�RI��W�P�mt�)-|e��g��S�A?���-���NFf�z�ީ���l�ǁ$��(�W�~�D�-�dA A�Gc9X�(ȓ�x��ɭb	M�i_�{CU�[�D�yR
�^ڮ����hnb	�#X�( �҉�e�Z/�����������2W"�F`+F��5	��W�C�f���4�Kz��Fp�.��dE^9�z�`��$�9	r����;FǃN�(��?�e��� �-	�T��ND�l�?�G#��04 �@�����|��:=����a�Ti議�vr����m�����}���|f�fcHC�����{�w�H���|��s"�%����{h;��jX`���e�4z�F��R��3�݈���<.F�'����2�.�4K��H ������:J~8�H��;VƮ�nہ�d��i�M��ϱ�'�9�@��d���j�������촆ΊU`�SXX{�[u����g�V�B���͹WU�)M`(��) W���F���� ����$|qe�t��Yc��>�'Qt�BИ(���Tʞ�w汚���t��(O	gJ��FW\����ey���v
卸�O7�r��%������b���z#��沫0��o��M%_kځ�sm��l�.=���o��?x��8��q�)��O��E��<Շ+�4� ���`���MDJ����G@� ���'���k%�`�*��r��*a ��ȼ��q�(<�H&�.:?I5����-B�,����� ��$��p�!�ݝc���*&�C�=���Χtu��T�x̕��6����X!�(/�*�C���y�6w�f�<�u&��B��t��3"�@M��y��{�E`߷K+�� �ݝ��{�hyB�	�j��YV|�� H����� ��,q�l�vcq�ӂ�h���-/��%����$B��7Xs��Vo������C��{	�1��0�ŏ!{�zCg�Q�K��=2=�@����(N���
�3IAh��s�s}��}����y�١k�ܣ�3�6�2n�|�#�B��)� ��sHN㪱��/�pa���M�ov�2|m�(�ݨ|���x��-8����#��x���Z�ʭM�v�L~�zP�6�+��Ag�|���+�Slԑ-��vVsrH�����6��p���H���k�:��b��v��3�_�Í�(������wZ~/I^���̖�IJ}3���˃mI����I1ث� erx�%�rEg�O�^�O"q�V�E��ע�Cl�J�z�J��_j/!�� ��m�Q�x�c�Ed��g�-a4��Z\����
^/�-�:j��[��F{�w�F��e�\���O_��D�����J��D�K ��%�uB���#{҈�48�6�E����B$#�������:�MK�]��~�q9Q�e` �>ְa��v�ǒ�j	F�:��2�f6l�@T��CErq^`��T���(����vD�G���{S���_T�"��A�-���Fkje��n�\Q'5ŀ��3����>���FH>��X���Pv���_͓':��&n�S���3����EGW�{M�K�n#���h`S0j�Pgᇼ��*�9e%S"'֐{��_`������
2r��Y�ɦᵥd�fq ,�19nZ0��o�%�fIh�d��ȡK>�|!x�h�8����܉��GC��J��bj�vH�v]xC<հ��T���fȅ��Pt��g;���c��jk��[1�F=+��B�?KK��x�D��Oz���Ե���u�o�J�9�C�-I_��J�3�^�hB�G.Y�P-=
+�7��$�b<Uo��qn�wb_��R<&���p�8e�p�&�����/�X�DٹLR>x5�:	�|���QW]5@����jw@7+#c1���\e<Y�rXY#N�%ݫAIgrs�M��ٛhu\�0���6�-��h�Fh�	4�SM�m���9�B��WB���(\b�	�Ab��w{<�a�ش�ps �i��]a!��a��z����I�>i8��E8k��Gi�Tq���2����\ϩld+ʑ��QD�>J+�U����M51�HV1;�{Č���J��՘V��^t�M(�5��G��Ò��U؊��U�-jKH�~z%�XZʔVu�=,"7x���q��+��?�&�(L��(^��S^�4�� �uɔ'gtQ�A�r�xK^ũS�xܣ��D�B����mi3��6��7�%<B�|��Z˟��]�H?LN%�/��{�ۺ٫OI��͐�p�`�p����y�JWQW�Y՚X��k��/�ݏ@\���*S 袊R���I�� ��Khʼ�PD�UųZ����"$�'s�R�0M,���?Ȭ�׀�xK5�}�"� 9g����&����2NoDq/P@�^�ԺK���$��=NCd�����&�Mf�l�g%�s��V�Ru�|��:s/�Ҫ��u=*AH�D����s��ӑ�I@af�`�Sh2D�8�|�y��2$�(I�ߵ�����nq�G��i�e
�x���7�}nr�S��Q �:"0s���n4�t=f���E��y�P��>Ow���5 ����V�_$����t�^i���\�����j�y�zId����E/L<oO�O�������8���R��>����D����+��4��Byf�1{��@5����3	�Fm�:����&`�����	�<k)�YKzߗl�I�;��>�ǡ���_B:ǻ�p%�8��e�z�����œ�kC�bY�8��!��u��f��j���Xy]��>_�l��^��
zdse5���*^��\�M�G��\B	U�S�-`h���c��\_6�5s) �ǉ����sPڹ-���.Հ/ɨї*,D�1�b�v��-������Ό�DEU�:�쳒%��W�tm����W�o4����|i*>v0<@e�j0l��}����R�妼l b�ʪ̏�;dN	�����3����V�a��a�"�A�����(��Bt�%*��c � ��L��۴=�P<Z
k�<���g�j
�5O�{!NB��4�i�c@(�I��E��xu�h���f��L��
4��@g(,X���*�{Ɔ��,l}�~�$�bN��6��68TFY#�`_�i-����{u6���7����9�`�Y;R�ˤ	�@��@F��q��2e��V}3X~c5�zK�*����8��YԦ�5�y�堆#�J��7}����Y�����"�P�TC�}`cE�ğ��	������o�zK�b}��3C�Е;{�^N�A��[!%ӛ]�0�D����ف@>_�/;?�V|W���*��E��)>r��?ǀƙ�1Vq����aU/A�<Z�p�3��1g�X�u��"n��3��y���r�C�u���4���N��9f��Y��p���Ic��C������5b�bmADk�3�2���H�yѝ��5J�^��l	��)l��FWaf�������~����͗8���O��ٚ9gu��|�����e���g�hGBt�[��1��qͰa(ݨ[�.����[W���[!Q�/,�P�n�<�ǭ&����Q��-BR��� tX��og�w�_b��#�rU�:���/�]{E��$�[z���bf�����A�5��aV�u��Qg�`R6\��Rx���1���rG��3Ƣ$wn����w�[�䖨����J�?*�(�85$�;���t����<�t:���S��d7V�R�@а^ё=���7	vo��]��#�~;�ZԖ��K�����q)�I���M~ as��#Ja�皩ɥRd�#nws��W0���9Q�3��J�.�cӧ�E��ڒwf���[ŭ�
h��3>�q&3lk�1m:��?�T�%��
�}�d"L��U2������4d�K���?��v���_��NH�έ�K�t��tGyT�o�WQ��L���O+�z���B����}f��{4�q��MA�;���[U���<}�wP�����)�\n�IB�J��m�-�5�l��XM�����g�b��+�M�-s|��� ��j������n+t=�oR�G�RY#)�s��˜��:.�dH�������75⒩CCP��5�Y��NXA+�O>�Q�i�X�Ős3ޚCH�}#0���EӚ���䊳�	B;#��T0��ߦ��e\�V�D�R�l�r�\���zj�C�R�� ���{��W梆!./�m���k���C\\�\iw�W��LR��e�{�V����ڰ���s�#�%��1�����;���P�� �.�e���y�7�%�h�Ov�#����z�g�f��c�g��N�ⷧ,�|�r�]�??�Y����)�B�m`>b7�x�����\ZяbxR�lh'K�`m�z�؜���gN�8j���:�%���^,��n@�:�$��� k;0�＀����qU���zJ���Z�,���f�E�ǻ��~��>އ2j�����Сzi�&�Y�R�A��M���iD/"!3S��fk7�/��_�]�8t����Z��z�
�C��	D3Uɩ�0I��PwL�z6P¤?h�xT� ��R~��[����
��#����p��ie$H�߄��0��{o�	��ݍo�h�f�Î�j���F�h�g��*��P"d��.���$��/�i�o��X6�����ARO��9���6���.�����m��|d;�+�Y�r���H������^���{F~�;}��_ڔ�=r��4n�2�P���r�?�jk���`���Zr�	C��1G�'�B����{h��Ʋ|��3�(�rS���p.Qv��ٓx�1xHn�k*�i)s��G�O�����qb�A*�jn��H�ʢ˸�P�st]�D�1�:/�Kڇ��/��8���s�%��4j��L�qV���D�K���5x�O����]�.�@qQ�X�"n�I�v������0�K��qۍ����Lz�2�_`<ӓH���^�Z�b�$��	�tK�]��u�r�D� b���-6���h�=p�Enϯ�:d]/�Ѭ&����T�ep�A\jp��}-���Z(f��pӕL����~��M��)4��J��N-l�4��6?a�$/��K��~�,�\>��?^�;�I"��+v]f��fv��F<9���?#ٞ�):4V���e�J ����C�DD!8��R
͜�W�8��;=�D��I�A9Ί�?�!���Q�����E�F<���+�� ��l��%;@Е�;�֞� �l�e$��}�b�s�F�"��A��Cš�m�r��7���;\
ײu�L�$��Ι�M�(=G��T��0����ಎ9� ΋������2��?ei�{��x� ��{�ȕh���HU���0jD�ݡ��������:�ŻDh����^̴�2�*[Mb�ej��5�}�;���e��h���L��=��8=;�W�7:��z���f���̹3*v�8�f�7'����q����zBBb[�b��iЭ>?8 :��/Oe�ר������?�XK����t���#��ǁ-�����#ǫ��l������o�`�$������L�����b�{-<j��y(mԃʘ;#��Z`C�T�Ϭ��WKs���c�o�E�>R [	Q8ɚL~>�l�Ғ��r��m�p����q���Ͻ���5�=��p0���qΘg���|6