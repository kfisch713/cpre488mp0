XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� ���`��Y��O�#�3|�l����#��,�>��ן��AP�����݃��V�2�W�}3q��v���k�'w��W��z�BjG�X"��Ք1����/���&����1x�n���]���dnV��y�����	Z}?d[F�e��`�a���`�%����Un�"�&��)��3IR�>"���I���n[���+��|�[-�t��p�z��JM	+ݻ�ŝ�Q�a;��� I�P#��ĝ�i�٩����������"Z��2HW`������B�S�l�G�IfG�EfGy<�$����Y/$�s�Y���c�70}��?�
iKҽ rB���=9��F��_�Ql�`{�a߄C@��h��7�ڗ�V��LtJв	����p����[�ѯ�y���nxu�H����'�tV�/�ѬC �]#ԑ-/�Oh����[��CB��<�<3�{yO�7]{4ϣN���C�!v`v���K�I�B��Z�����z�t��w�q�x�?��s�1ӿvh$	���c���N��~���>w9����?V,�?���?���x|@��W�.�:S2���I�����F0^�� �@���Nn'	G�IM���`ko5+Ҷ��{g���2K�Ȅ��&'��=R`��r�%a$����Pچ�.d��9�˹.u�"t�GSnO,�Q��f}x�>��ʱ�؂�i�LZ
9�d[9����4�i<ꭂ�۴�>�U�0�R����h���XlxVHYEB    dd8f    2160���[YQ�p��Oy^N�o�6{H�a~Y�u�4�|u�!��%ˑ��5�E��|�?5��ة%�iX'�zu�x+>�G1��sz�F&em�����F�������!&{��h���Is�����U�Ch��\�W�΁��e��ۭ���D���M��
��U��aH��H3��+Ζ;�}�]����;�6᫛5s����_����»��/�P_��;�k���D���5J^7�\2/��k�#����������� |/�/e�l	���%8[��3<���j���ؤ��Vx��u�ڱ��Yh��Ǒq��d�9�L׽(NZ���L��J6�9e���>�F�)��O�XM�rLd�b�P�P�Q�a�.YL��/��G~�-� +l?Mh!��L������{N��w�C��?�vG���S�D��9Ԅ�O�ܞL8B&�şG�E��Z*��Zqu�A�w��2'�8"O$4����}��x����_Ln�`I��e]4C��3r�N�4T�C9X����;��E H�w ѡ�e���z�޾e4�!3��T�ǧ�k]m��0���D��?I��D׶d;I�'�kk���#�zna��k��X��!w��aK�uP!��x5���1����1-`
�K��q���-�h�S{GK����[4iJ��uAv���tD��scg��A��\�Z���U�[[�~�8ה�O���� �8�y�:��uK�ƴ)���f�0�E
������ʱ���u�᷎����
p0B��h�Ƿ�V�Z5�ǡ�wƇ/9~S��\��@�L��.&��(R��<� �^>m_�9Sv��R	LJ�]��Ƅ.8~˿j�A�(z��Q	k�D�y�p�Cа����)�C�TG��Ok�6���H(�������z �*�&7�j��K���y�9-A1�	��fτ�]�%��:Q�|o��Mu|V~� �	�;e��@,�A�^�1*8�n@pw=<�#6���R�/O�߻���x"�i^-�W/�o]�ȷH�%���5�lLB�'t����3(�\<4נR��,c*3�k8ɩޮ�N��t�1a=.
����g\LKy�ᐴ�m�Ě_��H�q�:[�#"[�U�Z���?���-~C�H����ڀ�Qo@�/�"@��v����[�zM| �a�au0�>ǘ%P���x%�>7���#t�o���s������*��#��`j��G0 ���O�2��&���y�ָ3����'Ӗ�b�I����NPi��Z<��d빙���|W�%w�AS�pX�<�^���:�O¦Է#���j��5�_�e��Y��=\m��9�T,G���E�{ڜ�-�����QX2�'M�!ۛ.�h���J����
��b���ӯ�~k��������z��98�Q|��z��;l��w��v����87�ZR&�E>b�^l��+��$_�&�Q�o�Ȅ��t�[zm�0Q�|��e?����L����ߟ�3Fp!�jW�����s}�	 ��6:a�~��e�U��%Ғ��=cp�lMX������R����[��G��	���1?�7j����hq�53HV���T>o���R�ߟ{��B s�S��Rz��@x4+���u������==��`6\�2�ۃ�W��<�ݨ�j��te�����U���5�.�}z��"t����m��Df����#ā!�5q[Ť^��r^F����Rl�qǾ��8G^�ȱ��ux3����\#Ώ��{(&�����U�>aɳ�_�<��g��V����"#Z�˃��q��Do���� ��{�Ւf(#�qWJK���>q�9�-^{�a�Y8����1.�z�m��h��p�O��OqcDc{�9ۻ
��Z�tvd�$�{@64�y?�T�;'��D�ԳH��g7��b�t�EC���sr
<s.==��u�m_N��
8P��{�Z�|�c2��ccr��څ�ye�ڹ|#vQ)����)U<�/��T�|:�fj���6U�H8qf��X���߆�π�N]��5��J
�AX��V�4g���r=QG`&��]�k�%�!�'9���\��_1^��X�����d��h��ē�bs#�=;�u��c�!^h�;9�}�t��M���#�}#��%�
L�4�'�mۏ�Q��I�A��2�<q���!C�J
n�DDMWZ��*��+�}`6�K�>0م��>�9a�=O�����#_������px�}d��2O�� ����<�(��b��L]]�MX���@�'���I\2)�B��K7/�M|�gG�q�g�I>����Iʅ�fH���O����*vl`�����k菺5�u�M����s\��d��[���*lo�
'�4N�˳@,r���Zc��ms56���F|�OE�p�L#�d u����1^-k�n��KW��w���Q*��|h`�&lb�+F~<�^�����z������io�o�c
R�ρmA��b�Ȝ9�,�P*�j�^:��E��qvB���K\Gt5��=�G)�'���(C`�:�4&4��|����5��:�~���ML�j�v�kt"�]�n�W-M�_��Ϭ�/A��l���g� ��C��C~���4���������SHp��B�ɯ^��ʠ����sٮ�W�xj���ori$�@��h����d[��@D�$No`�N�)g�lQ�ɯ�����"{��0���P�&��� �������@
��>��B>x���"��'�����.Mo�eo�1����q�D]�o�o%C@����Q;��Dפ�P��r���MiHU�!(�"t}��'��V����¶F�K��VɄ�UnC���7�:+(ւ�vOl��������@�H�[�=���vۗ@�|�]nh,bإ`�w�I����8س��Op�Q[�Nc[f�UR��9`�d�{�zbs�"��_V�aX�f�cR*Y'$k<�I1�t���F)+nrm�0}F���
��V��Ÿ��q��b͝�s+�Kp=�n�`Tf�%0�
�2�Ub\=���r�Յy�e��az�5��v?��`��MPE�;?����w�?ϖס^��o���o�X��0�#nD�O��6*Ʋw)�����t���o��V��_s?!1a�hC�`���,����B�`:�,\@k6�5!e�>�fP4�`=��s�":-I=uٕ=u��8dޤ�C�%�ѓ�S��>��,����Y�'�Ͻ��K;ܨ�yh���w0w�!�	���PR'Q�~X�!��C��S-8�ˏR�TN�<�i{�ѫ�*��(��n/���ix�+k3��4-�]��L�r�ڇ;ƽ{)A ��]�>�2AM��^4��&�N�Z�R�j�ГR�I��M����_�B���ڄutV��q8�+P|�g�fc}�7��a�{7I�`ܟ{|�����*4(�~@� %=�Z�_Q6����H���zh%�"9}�6MN"��)(��P����<;;t�-GV��6��F����cko�CFqi쀘by�����- � ��'�N�fۈ�m����^�6_�6���=+}\�z��oi9"��IVY�'�]��y�[
+��M��p<
@WEx1��4�VpbH��Evjb��1����-iF�d��Km�P�Ur�)tW���w�˸x�*5X��L���a�Yazi���Q����<��ɏ�{�G*�(�RMi��n��D^'��;�1ARos�,Q;�t/��N��1��v9��̾.dK�<Yk�Nn1��s�꛶���~����A�/�J)I$GTL��n}L�/m�;wU���:/�<v�S4��զu��勼��~:N�X���$/���~O�ޙ����p�i�xR��@��Q#Y"�?U������m��B�j8�  �P�\��h�<�? �<��$,���{�0��2�}�{��*� ��� (g]��\2�zv)��@ULD5}���\�YWZ\.��.�y(,�^fI��Y�)��g~�������u��j|&S1Tj���D�RT�;��|�X~Y��L�5Ƣ?�?nud��nB��m�/a�Qv�:7Fk�O�$\@v_ǣ���4��V�TT����w���5zG�;��R�������k�G^ �K-�	�nl�?#��F�ɼT��.N����K�1l1�ּ��ڛU7��p.#����[h���TA��[� M����m~���%f�L���t�:_����fYk�i���c �i2GȽu�������+��u�-�܀5Y8�FG���Qf���ЃI�%��4ό�����a4��w�<�k-[��e�T~�h�]����!H��0(t�+�ވKVtL�Y����{%��7"L<�s��\zI~�ܼ�ts��ט+�!�>4)�6�g���"_Y��S���EL`�f�������UQ:	 I��~V`2'�XWGo\V����bJ��X �����oa�L_{��r���"H���)"�1�_f��!��@�;�5��q�"0�$��'� ��D��V�M<���M��`"�Q�(��bJ���E�[2W�Azp�'�W��´d�ɉB��-	�?�GBV��#T�$C{��+ӆx�5�ڠ�rժ�8�_�9��T���7IT�J��&��ɧ]��w�J��=��?�/B���䫱a���������wz ����@�w���)�*�PBeG��%�Y���o����<ql�$�Iu'gN� �s��"�`8�T�[��,�dnu�_���E������#�l����n9�����tP��� TH�*뵚{Cu�P�0��E�x���zZ���J�7�O���w9� �ڀ
��F�[�� ��k��9���p+=��nD��h7����>�P�@�+�L��׮6�&���	��nc���n�'��)���m����hs{���/���^S [#���ſ{��t�*��|�m�4)>2I�'G`�mcN����B�^JE��}�t�_:�������0q>�T����H��o* Пͨ'��_5s���-Nt�����f��u2�~��5��n�?T�B��p�͔��D��5p��Lّ�T��Աk��?
d��C�hO�����y^��f�S��<'���c��_4t {#x�p�Y[��~�X4�y��"�78��;
��@̭;*�@U��j�r^A׋����:nbԨd�f�~���O
�sYD�їUl�!&p:6�ۘ:Iu'	����'
�{��szW{��D.�n���֑]87 �S��v�H~R��� éɭ���A�����m�`f4!�w	����?�Q�W���g�Fs�Jnj�A ���.�	k�JӒ;~J��Z�;���mmм��'	��%�3@m���ޅ��tD]��(�����w�r[�<M�1(���T����4�\��ƅ4���b���>ע#:�S��)�X���d��Q��~y�Z��Q�6&���#�o�#����X6�5�^�sZ ��vu"8�xAN,�Ş����G��!A$Sw�9&ɽc�����
X����Dӄ�$�+�)��>B)��p;[�	�Y��9�R��7��|��!��(4O� �c���(���.c�/7�6���/L�Vajfz������d�2��$�p��Q�bHI��/���+f�TkA�_�]��xR��+��Y,o�~�����P��v�.����f��v����(�@�Ȳ6��f�H޷�4�#���/vݛ���ңt�����<S�S
��l�݃qǯ�4�7��^i��nu�b�{d)���
��F��LG���H`�W���@�YI�D���������Jp�
{jY�τ��ݦ.��"��@r�|7e�,�m�`�%/��Xs~<8$טߣ����� ۋ<ىmX׎����U�F�3��az�d��:"�>
����8��c�X@� #��X����yD-\�f�=�c|���{̪x��P֩�� #3�Q��RL���o{�4��	��1�ȯ�]��)�U�8m�C��/L ,���)�\�,A/�����c��|])�l�1�BDw��
z��;PS*��S�'�y��iv���R�pg�R�EVh�Fҭ�\��<r|D�ɒ�ʛ��w=��6�{�j�X6�>8�-��Z	�����{)wY�\Y��}����5S�H5:�7,�Q��1ip)�J��M�M�v&"t*���=����Č;z<1�jX'��`#��
�.��b����D�H��sP&����t���L���L7��킲(K��"�'��V��%�>�K;˅M�^�J�8���B�q]G,�(�A�u啿����\F�Rr��� B���T���9s���q7�^�hPG���]���Ql:� /.ǉ���Y�R���K"ҙ4�[4��W.DY�&���&�Ė>��M,��a���b��$z��:�d"sb�8�ٛ(�}Р�l@(l���6|�K��BISu��@��P��m#�&Vɓ�W���(�j0|s�M�_����"����L
���>/a�Ŭy�{0���������Tm-q3��×�<��$�|xm	c4��yC��*�
/	��#H����ԍ`�	��%�5����1�W��s�H��oy����C!e�z|*�����j�H�
�j�o�u:�E	Rc?�S�-z%]�w��z���g`ߖҎG���l�ɒ�PKx��6Hܚ�ȢE��S�ς�U�O��R[�2��L\GI�G����|(��d��JtH� ��+|;���ma$������**�6�P���[R�W��a�� �xDS��/6qΈ�{N^	s�����1��~��|�Gou6�q���OݟF�̔H:;(��yt�`m���A7����&��B�f�VI�t?�d�C��?������wt���ޢ�FB
����p�G7��X| ��j<�4�(΃�W#��j��Oa��`J�����]<���]P=�˼�����)|BI)d{~!~�z�DvK�J�I&�~�9x�C[ ��(騪�u-l��YR!�j����FI�e�"a�p�~l]��mN*D��-��L
�S�Ke�!�"E�w��l�/N��'DW�42��#k2��ć}��OE��*l��:s"י���`O0[���L�"�KT�zRj��� ��i
�W�J�$2��l���=��|��@d ����\��o�'�Ԇz��0��i�*��&ݰי�_Y/�|�k�Q������>� e1����0/�&�� \��q1�(KD���@h����sW���"}�q�k�C
���uoD��^#9�����r(,� h����r�{;#��H:O�l'��9�#��ٴ�Af�D�/�]
8�*�@ܔD�)�����rA�5���Ɉ��������jg\ɩ��@cǞp�	���������-��|���JVy��0��h�H[N��K5�x�N�
�Nc߮c��럈�x�v��F���E8���d�K~�~5����y�Rn�5?�٫nܥ>(�\{��pX�=�Z��zun:��I�o��z,�ĲGl��3U�H0���m0���2���Oa�3�&7�SP����������J1�Ey�V�Q���K���	fꑖY^k�#�^Vc[�m.�H$�?�S�nmy/��r֞=�K�n ��`���tO��5	1���N�<�) W�2���ҏKa��],�FV�<q�1���W��[�FA.�J<G.�������t3�h������������ ~<��%������a�J�]<�Z�YE� ��L��~��&:hgY1�$��*���%�n͡UX��wG�������(��x� ��a��grY�2gѠ[g�c���U�A���l1	Q3�G֏q�^{��j�Mq����RS����	.�;�������S�2c{�z5�gx8�n�p&4�8�57ǽ@��i�I�����DqH���ey?�c-�jQ	�dUf�NLΜ�S�tB}ޫSBzv1�FlG*h>�z;��ny�e��o୴Sq9��t���TTZ��J�����;�d�yn����/�Mz,xP�[ �#�p0�_Pڧ����	��T h�F��8ڿ<b����]B*�{*ܠ���z��p#�u%�F����X� 8-�<�j��XI�}!2(���U$�7�D�+��3�VJ���"e�/ػ�Q#��=�Wo���XQ6��I$p��BE�o�[kVBV�A�XV��}�.�R�涆������قu��=����_�$�늭Y!C�"y���F���F�x<[0�91PV� �<z_$�]�+���;DdK����=?�˹�}�~�fH[e���$��dSlLa��D1g�9P<�X�
&6�3U(�~w�2�d�҇��va~%���fS��e��;��r�pǝ`9�~��ec�;S�H�k��Nb* {	��}�}��\�'\��m�h�z����B=��y�n�@fh���B�@IR�X%�������#K��