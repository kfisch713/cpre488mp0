XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ٍE�\<Wl�C��M��80�1'[9�>:��+f������V�]03���ǫ���\��,"� �=� �Թ鋂����<��lz�.�c���t�P41�>��}Ѫ���ӊ�&�uz���v����5����Wc���ه�wc��A_�Yxr���w/�q��t�
���iC�W  &Sj`��h������S�;�3v�����t �}�Ϊ�3���ą�GN<�o�,"�6_�IN> 7`/�iKz9�	o�5I2�R��|X�a�L��Vmh�/�v�_�����a� nl8�,��=??�z؄�&S�m&�σ����Utbv���?�K=E��ֽipd��X�ȋ����_u�U��c�HO��Y)�;%�dc�2Թ�D�+���)�.��_�|7��rOA���� ^2S�wS�
�vѧ|�y��@��G
��)f��Iby8l��gŞ<;�
Ã����pU�R�V#,T9��LG�SԧZ�Ȗm鮯�_�o�e�&o�*�B�6{&��6VN�n��G%��	�f�Ʉ��#���4�-�ͧ]� @:�%��R���8�G�Q)'��k �5QP��Ă �]�\�/��]p�NAM�B��t0c)���#<ps&����y1(ģ8�P��v��� ��W�+e=Zs�K~�+R)8fi�?$�D�	P��[tIA(*�Vg�fs��K$�l՛���M�D��)l���h��8��Y�s�oQ���>���>^���F:����x�XO�yK�)��"�6XlxVHYEB    b3c6    25b0?ҳ�\� �q���w ��M�[���|�'���r�g���p�a�m]+�q:hB��&��I��r��L�p�w8��K,`�T}�.��`I8 y�}&����Q�@h��,�2�i.:�A?Z�jV���F��;1d1�7=a��R���?J��O���Xi#���aM���=)犡7Fe�����W����ƣ�_�������89�;A1�r��nNF����T�5W�Q���+���2v��rૉ��廔�d|����"�ߊ;�r�I�z�U�I.��4���	�U���|<l�4���ܰj�ܫ�|6J�1Y$�F��v�$��/�5k��pٌ��0��~x��_���O�R�NN�G)������L��L��<B�S�T%�ռ款$bG�lك���#�uT�j}~��(N��zz�=�A�J���j�j�D���1�����9ӊ�v�D?�/���=���Ff v�:����T��o�f�c����00Z]��7��������B�U�_It��>������.������aѧ0eyRD_�i�ֆm\�����	ߐ6%���;�C�x���6¿�&�sᴲO?�޾�0r&ɸ�w/�c[)İR�A� ��t��&�p�ɀ��Ln�s�0��'�O�]���6�i�諓'1��M� �P�:V���p;�\���t4"����+�5t0��n�:�mI�����b)Bw˂�]	�U���X�=$ì��p���8�2�4y���7-4ɣ%��j����x�&y�nL[����,A=�ӧk`Y��S~�K���W��zY'-c�폻�9�!Bl��i)���A�jH�Y|&#/�|��O�[xo2v���Q�,[6�j)�n�l�i�"��ݙ?�h4��N��{��[-�* m�y��)ִ�lȈȢ&�Q+�sW|w�`�TԞ�V@��x�B3+u���b�E��wy���!�fT�ej��s�7��S���57:5��o�j�f5A��D�H�w���]�^� ����'w��å=á莅�9$^^�i���������tN,�8��
Ӕ�<rF��d{�2'��1�gE��s����yap�.˝,)�(�ڇ�;�.Ą�V��T��~C7�K'�t?>[���}@x�<���J�㖒����O��L�����@�<߫��W7T�K��'��i��.}�.)��-z��6�/]n�_�zkc?���j%��ǫe�K����K������#���� k&�S1�V�������t�-W���k}c�����屍�iHL��-��ژ�j����G��φ�XcPm����Dm����ນ`���ښU�v�6��Ů*��ɨ��{���d������
�t�5� �\�|��YK��@��e�����S�7�_�Hn��l�>l^�+����~����0�].��4X�gTO4<7pK �l� 3"o�Ů�?��Ijp�Ÿ-n�,e)a\��ƍʒ7��Q�1�R�R���Ѹ������ރ�Ryv���� �}a����}+�0U}����U2�?��.h��BB(�ĜK�Bia���΀w9��gB���L�}F8O�����n�k�P1���zJ��2�,���yK8 ��-��I�^c�?�Y�TN�B�u�+�Ah�K�A0�42��"$��c����(�̟�Q	v��p׆��=.��l�9����f��av��X7!H%uS��f#��)��V$A��+�R͠|(5D$����a�i@~�������~�oA�	f�/�>7NKGIg�R.��C��Oں 5�ʊ	$��^��iu:�	�e���g�z\4��o௦E7[�ٌDBy��Xxɔɋ�'�Y��T�$�?,�u�(�/��4���㪑�U@���!_��E����MX���X��?2eyb?��OS�r:�	�AK~㮿�glV�-�ʠ�LΙ}ի�z��Z��
���s/L�z�H~�ɜ5��ρ)�~���;�+�$�ԗM���-�]���hߦ�#�>c���P7�)�����	���p���5����5Wj�W
`c��@�g��7�$��N��gX�T^� �ת�=�8�$Y7��b���҄�S[���'35�2lZ�UYMӶ8��ۧ�|�6i��C�14�V�#;�[Q�,������,vE0���b�u���hd&�'����e}I���Zm���ۘ�6���O�f����62�N�����&NNQ����T����/^B�h+
�?��M�p�;A��bE��F�11>��*@,������j�t�F��i��J����Թ��N����k>/��w���e���i(o��������N���>�F�z�	�g�f�v���	Fj���s&Ex���c�!�V׮^���&���}i����u5���W���P��+pOǆ>���·� T�a���&U���YW�*�tl�I?��L/�M��l2sC�,ts"-����?:1��T:*�8[>�m�h<J�Z�����e�Z����y{�A�XR��v�`Q.������75׽�S��4=��=\z�e[��5�qk�Ne]�:�ٱq[��cv���J�ظڑ�Ȕ� ΐW�[0�C)�� 6k� ��1׍���G���L)�ލ1a" y���Û�\�#����umcrh���O�ޘD��D�<V��<�$T�(�%�VtM�z8�B��C�ha�}F���#/� W>X���y�DrT��rp�?ɸ�oȧ�_�S��ʋ����bH�#��X��j��ⶍ�Npic�����7y��s�N�Ng5��dN�ԲpO��u	d�	�G�^.�,h�,�����6�iJ�"��`�s��@�
N�픔���ժCRs�.9��\��a9oMٹ��Y��eh/#�)�$�!����k��=~��ըjؽ;F�f���#�԰��G$������9�I��UVϱ3��T����~��3�r1��M�E�4��[�0S��Nn ��
�R�4W���?-u�A�uz�Ҽ����]�'�ÿ�I�PCa�&$�錉k�w�FiOM�+^�s��,��L�U��3�����-�Vr))�U�:���B�]
3��Q��E9�1,À{;���+�7�@��oEM}W��_G�&��5���#�i��%�VQh��۞��ؒ��}�I=�)�M�cwΓ_\�%�7��]�O8�l:�<Ӓ�ӹ~���P�7[��=�:уQUv^B�Ѕ=	D��i
{=�t�̛Yv�;x��b����u��1t�e ��V�o94$WL���u��~@A����τ�7�U�t�y���:�g!��Ζ���.��� �������1�{y�X�3�ϙlH���O3Y$�A�؇��5?�����	���s������Q���
(OB��%���r���8 �F�����a������&3�,=���6������1��R��
!I0�wf��i��`���U,������Yv����p7�*ܬ�����;�Q�ң۠�R�$(Q�>S���O�6�����q�!�ka!������t5��5�qM�>t�lq���)q��j��/�G����0�X�����~��^3�O���[�	�6��aM�g�ÿf5Y"�ȕ�������5�:����v�	����'m���I�=bw A"����"]��j� �QC��jnX�mzP�����^��­�w�",]5��W�{�^�8�(�(���sc�9�|��7D��I�����8��r���� +�г�T��O��d��	8�,���Y#����3�
(��@��J��sf֞��֯p�cT�o�oo��N��i)Ml��y��C}��<�ǂ���Ǘma�5'9Fx\�Fۀ�I�U5ŏ!���Dt���٦�����z�aڋW���%��y�5BArEVX5>5�X���'���i
-��~��0�M���@�[s?R�������v�q�� ^��r������N�6#��y�T�!�JT"��QRqV��V<�sN "H��^��]�`J	��3~��l̤�
�,#n� ���)+�'E��~�bd�� Jr�I����釚R���Ճ=��N1h?�עCӈ���V�:��$��ڳ�]O����������(�t�=�MwXq�{?נ�������N�?e�S�8��s� 3ν���7̡�\�/�X�ĄpZ$�sX��YD��v��9���8��픨��kU�$E-2�����y�4)��h����;����{գÛ}�H���P��@�5>�>o�c�|5��i���8L�5�2��>AϮ�_X`���Y%�Xh�^�:[�6D[r��L_�/�e���O��4�6� �q��6U�K_�ZǊp�h-�}Kt�o��-�'��9\ŕ�U��E��6���Ss#��Ǯ��8��=�q�ڎ۱e���m��~�۾��:7�7qr[ip�~w�ų���|���'X'����ro�{�I���ػ)G�oǟP�[|HV	�CC��
���t/�k3�ȏw&aT6�v[���A7�#k�/�N��y���}�$�Q�;)3!qk�מ�s�E%~���3p�7=E�kŒG�<�w!պ�w�� E��싿�cB*Ns�
�E�:��`��W�R��^E#e�=<RY�� ^n���Q����v�!U���䂱2p��ݡˮ�J4�=턴���n�`���ήf�#�I�?3҂Cxʢ�W�^b�p5$�V��rP��dR~�bd��q��Y/D30TS��_�c��&��ʐ=k#oy:����15��:0ÏGb��	���]5����*��Iя���d�u�%��(P|I�����+n�c!� ,1�
�O��+C)֋��K�دÑ�����m��n����]~	��E��Du�L]��Œ�ϝ��î�ͭ�-��Di��E�WWI��6��YwFL�(�n-�ƹ���52}�]��II�K�5n%5�"�(�)���Ҩ+�m�δ�fD������)�p<=%����q��u��촛bD���wwT��)�5�:L^������}=�L0�"ｆ�e�Q�u"�01XV	ֱ�<�̠=�fe{�Y�Nxk�����Z���O�T�&cQ�F|��{�u��SB@t�n7̳�Z���+�0Ȉ:��j%��䕪h�����D�a�N��Y8�Ҥ��u�!ڱy$�C����{�B�	אH[f᦬�V	Ɇ��u���AWG/Ueh�`�1]�$�F�y��淪�����G�F(4I/��Y��.ʣ����T��QO��e �!�.�6��[.����-��{#(ߠ��C��#Y-,��L��<2����5^vK�`��~/��X��K<,��1�y���K�*7ҍ�H���X����-�ѻC�~K�
����ם1[~%H����ђ�40�ݍ�;;�H3�xڜ8���N��8{FZ2Y�C���O�V��Tsz�>ک�gSf���'&����e��2U)R�KW5q�<*�)8B�(�*UC�Ja����ǲ��ֆb�Ɋ+S� �&M�\�'�6�>���c5�&3��n�p_�[�&9�n��g|*�F��q���p���f3Ozh���&�g�����8�^!z��ح#m�X?��&]�ڟ^�{�k()U)AW4��! R��f�F����=���z���^5���K��~L�D�k�'j���J��i�+]�L���HW@�� �#u|���}{����HX���\��xX�5t�����O�jd�-';���$��L���+�0�����T/:Y�Z�}��9_�~�&�F��EpP��U ���mb��箤[���"=(�S��?D�qS*�c���NȪ��ě���0]����"C�8�
�(�m�J{早�=����}#���fE7A�j���ͼ�(z'���U�.ة��b�S�g}&�a�!�[5K��O�W,f��[�)�F �&J�%U���9�zl��V��eG�,���e�u|�m(+۸��6�҆��������a-z8'��٪ǤiR�5&X6C��c_v�*

#��/�f\r�=t& ֱK��]H���^u���E߽�:I���Z��rP���<���T\I*z���h+�U�l�Qm- �@���#'1ʬ��ڛ`���@`��D���I��A'���ΔN�|�7�w.E�Mwb�fAM����(|\6�9�,��퐭P�G8�0u�ֳ\� �B������!r�IX��ϔ�{��=dy��}ĽM�Ѓ(�T_�z�9`Ͱ^�Z�p�G��$��o���=9>��2��ޏiseC/z��N{�f�Z�:�*�y���hnG�.�]��VPE�aS���>����O_8,W2��?fO�]��gOn�J#١#)��$������\��� ���͈��'�@a�^(6qU�l}�C��j
`�H!M���ˬ7'vaL��Ԉ<��*�*"	��@:�?��p�#_z��r�Tx%i��,~�Vix�M0������]�C��_���{@d�jww��	,st�ߛ�Sm"�,Ϫ�\�&�Md� �XzB �1������ x��a�zJ�e��o��r	À��	{�x�L��Hf��-����1C�lF|�K����bRJ��b,
���W���Vl�ԴoNSĞ�*��M���)�(�׋[Ǎ��Dbɛ!@�Y_��X�7
������Ţ��EN%H}Pc��$�������N@U��#�3_��,�:"iR��Rj��fz��A�P���B���v*�0�\��"t��l�u9-�~j��t�Ѳ�7ҢH+r��۷������	���Ȣ�@X��(.�0�RWb8H�4�
>�z�GR��0��ތ|9�2R� 8�z����P������.��n�X��~H<z��I�e�6�S|��7 �db�]�R��8FF�USˌVl:���#��b��y+�H��~�Z�^������9Q��s�h:�	���)8'���4������e�L������M4��뿣3�4[��͞���(��";'�2�G|8"���t'w%z�U/'���:�`����VŔ�J�g7�Ѭ�s��Vg}pD�Q���/W�y�o� -�Y(�@�x�|��ӝr.����'~1�r��v�d�r�\OI���a�o(�Д2��^�8 TE�p�k���/G峍v�@�*(���|&v:%4�v33^Jw�g�-�ʗ�켻щxf�%i�Lٞ���V��������v�y�@gX�������4��G� t�))�y>5{\!���w3 v����t���7R߃Hǟ�X��`�H��@l�����ZˀE6�/$h�&�h�a��o�he�/f����l}@9.lŰ�7g�P�DQ[�^^j�Y�y֙�R��(�ݔ�������=�jd�t�+uH�H����&%�8��	*���耿�>�۝����9����H��H=FoR&
r�iFI𫚜.�"�z���7_�*� ~�L�01}Cx�������x2K-��ў�G)K=ӷ������,˨�W�d�r��
���(e5��= ��{U�]���'�1��ϔ�rZ����3�Ϊ/W�b��ݧ�k+1x��Q�E�	X�8 9�r�{���o�i�i��X���ʚ��u�+p���
1n�_�5Eq��۴-ۤ�̴ֳچn�v��5�Ɗ����Y�m�i����|s��-p������$r�źyZD���~�L�ِ�@m�vrs�FbB
U͇t���n�6�,6��q0�fKĀ���uj{�,���e֢@m�D�H�r���h�P��,�<HnߛCc�C} v�	>3{Y=����`_v)Y.��[���ߚ�Mk5]jX�~x�����'��粷uV|a� �±������r-w��i8b+RU�{��K�&�����Ĝ�o"��I�E�2���E�Q���y`j٠�y��Pc[n��n��f���H����1������,��E�]�Jj�hBS��8����:�����⨓�9T�l�\����W>��)\����u�|ڵy�TS��������0u��K�	�l�Ix�O^Zf��Lܐ��ޅ�K�ޚf�L�8����-�E��V*��t�ʠ��B�x;�$��O��ɶK'B��D�����_����d]P(=�-/��3�k/]���l��+�������E�$�kt]_��b�v�_lj%&�КT��`�h*��P<�0�Ԅ�[ >����d�_�7�1�-)����Gi+b��J���ۙ����=��K�y#�3ʗ旟`Qr��\Y�܌g-u�O܆�|=n�1��X�*R��M�~�<L1߀\���zo��U���k�Z�Lr�S���a�|�Sb>�܋m[;ʚ.�POOi3���a�Pb�QweA+�{bnb��H��5����$���5��=zF�J6u��1?O�э��F!B��QQp��M/�V�=w�S��6aM��P�&����)��w��!�a>�w3l��g��e�:�! gB���*M��H��=[l��};0BD�Z��c�:-�	UA��<\��*#����a�>O��!Ψ�T[6d�n�}T��1'�O�d�Ę3ݙ��?��s�Ti�I"�?�*���0_AL�Re��昑��j�>Q[����~EIh���F��!�`iK_���I6޶�Ǎ(& 9������j�nr ��@�ڱ��':xR�yT!{��j8�u�yB[� ��`�c�

?�+�1���=���R[�H�Ҍ���V�G�y�_ʲ� ���N�HW��GHl]���anU�mt2f��ō�P$�_}�!�����o�U�;�D#&��;��/y��RB�(�ʇ<��M��)C�ڲl�f��-�̦A�EaT�H�8y؆�o���孬����|h� ��ʆ�LA�>rbh�Z�m��Ϝ��z��*$�}F�K�?������?�ց�����PH�s'x�V�5?������Ip>
Y��܌�F����#��lw� M��8�$�&ۄ�mw�ı`o	]1�q:|4"4�ˈE>a �[�e�Ŏ�L�J�x>��_��REGI�*�� �'�-e�Je�7�9�=] �X���K���9�)��꺕׬�í�յЈC=[�*]�ӷHI���=q���"���Zm*eHȪ�2�JtV\Z���,�,�x ����xɥr��КF�'�-�(D��v#�H�~+`Kf��K[\ꏟ�_��=�g
}xN�PW�ꢵ�͊�
���y*��=c���6P��2>�Y�b�@6�վ�����
�?��i�M�U;x����pr����J��q�v_D1١�5��WJ��ű�̥�hC�b�ب�	�v��������&�9�����+��/�	�I�=��@�1ۇQ��O=��T0�O�CM|̓�M�����[�#��
A�鏹��2d^%n�)���"���H�j����>�Tdj��@�=����!�CՒ5 �^v� i��[<��)��^��7��1˃�l:��$?vW|͐N4E