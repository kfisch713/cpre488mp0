XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���%������0���:j�^M�b�n���Ap�U��:�Y��d)��/���fuC���M�k2J���'p졆0����y�����t�n �������bS��U�:�rr��C����q����`#��pXV>��rS�C�['����7���(:i�a�rIݿ��h�ý�H͉�m��׭TD�~M�	bL\�c�3.��oav�o��g5�fȄ�$x��*�����ԟ<�/�~�Z:�m4I��vF4i����c]�'U+z�p�
Vw��َ�k[�X�ƾ�mb�V�Rݷ$Ƹ����;b�A���t�ģ�ǔV4�T**�?��TK�Y��J�j.�����21�x���j+s�oԍ~�v_&@>4�8��J��D̀ {sRH�X�ftr���F���۪�<7й�|*�F?e9r@A������c,�NIY�o�q|���&��)r�_�}
� <,�/{���%��XgF���.��U��3+G�� #o�e�W�@�l�V�O,��i/%��F��3?�ghG�E�t��/�7#qz����r1���6T�	�4��Y��x�PȾ����p�Q/�e�qEm=Ph̀���]�-��b�h����L��21�����p�]cw���
TEiJz�>�6�U�Ol'�۩⚣�77��\t��&E^������~gak
����<*1�B.O�"=����	��� (���h���>.I�rY$>g�^4,k��P|������:{��(^�+�f'�D��XlxVHYEB    42ae    1110P���.��KHBZ�n��i��xw�/,"� ـs��� +�("�~����dUF=3�	
jR��O�Q/�'ZMapo>��h`��[�D�Iiv��(6|���
�6�ݧO����n�%�~���1����LOY�O1}��%HRLE�d�I�6h�a��N]�9�~�	i���V-�Z�>6���ٗSP����C+_�_`=8L�Wj�e�D��G�e���l�}�La�_�F�ׅu����߯��q/��!ȵ��
�����K������̈́( ��򨓵�8ү�d�5@���؇��<�N�$�p
e���'�R UmiH�e�rbfv��O0���S��4�_��=���c�(����g�1$�!�ٶ�A�>C��F�%�2���߰��g���B
�	�t���6��U���+���ϖ���i�H#4��/�+�͙�j������c��E������SϷ��M&/zr���S]$�M�4f�"���]E�0a�W���a��-O�=(c�b�.c
u4��MTԁ��"�²��o���^��ʞfӮ�R��i�ǍbVѽ��T��Te�Du��'���\.�
Q��
���Gu��`��Hɼɻ�-��s��ʵ�m��<_:�3����"�lw�@.�"
�z�	���<nxqG@�������]]�;�P�a�q�vU]d2����D>�8�1]'hN|�N��@��X
6ϊ�J��=6�@ �8ͧ�T���kaҚ����]���qZ�4nc������lT�IR
�f�D����E������#A�D�,���TU�cM$����0o-�� ��S~v�/o8�*�ntsu7�d����ڀ�q%��>Vǹ��W.WX#v�	Nn;T�M�b���
�\��*�eݴ���G"�G�W��u�O|��d��&��B���CY;��[����C��'K�x�?`�Ň�;��~���r��}�}�q��"�R����[��F�C,�n�[���JϤ��[���'&�֔xV��tZH!��1	d7b�L�}��D��^r��� 1����pn����>�>$�|�W��-�r�xZ��}�Έ�u�B#,�	�kƵ��:��V��~`�t"^�����6���0kt��`lI� ��8����O���Vm���� �,.�4��q�I"�樂0�3t#���0@��s~2����W{�Ɲ�۰p����{"���i�>�D�7.���Mb.���HgK"���mrGN��0f1���m~�!�f`�Č��k�-85�ə�����se7�J~� (��������}a,Yp��@�����^C_�A��y�d��0T<|�ƞr��7*%#r���Y}�� �;��՗i���؈�?%�_~�vH:9�tA;#мP:̆T\�*�h�����?BYu�?��E�O��W��q��H���a�c%����{5o0�vL�s�Y�P��
@.(��8}�E>U�N�4�2��A���GC���a�r�9�8��G��>�[p�j�w7e�Z����8PaK�!q�<9Wɹ}1�^unu�}��ڜ�a�ٵfGٲW)�%\;�#�w��e���eu D�Buᩐ�Qi��p�0X��S�D⓽0u�~Ȏ��)t'g?��q?w���L�%��ם�nY�S�{u�?���􀜏U�|��k�\�����h~@����{S��1v�#/�E~KJV��#)Yl�F�{E���Ʌ���![z�ߎ�汨oƓ@������l�3xh��5�^[��'f���EL M�c�.:����sʲ�d�K+���N��Q�;ir��:�'9��>[)k�b�\�`����]ep��Ď~H�tY�ͬ�nTC���b_B����� �O�õlM�̖
O�*�ر�q�!1v��e��H{2�����a�'N�'����?��*��|FE��ǣ�Z'�a@���)�`&p�ϡ�4�e�Am����ƙ9H�r�P5/����v�a�Tb����0�WK��\�n�	7�)�u���4@/�2o[��d���a�G�;	d�Q���0F��z�NN��|y��>�r���y[�̤�xx-��&N�H˽鑘���ŏԄVn6��^���X�8'��\ ])=���L0O�|LC#�k���U���츝K�C��:3r(���8o��`��j���m�U��Ĺ��͝��W1F2#֚�bc���.w<��#���å�Wح��e�юM�2��2G�3,�����Z���RQ�nCTғ��r�侏SG
�ox�}��E���£L?�ͮ���i�uA�<�ɹ��:9�'��?���a%����YeMa6ZU�5����UC��^�$H5u��Vܤ��ʃ�^�A���0�x��kn�Y�����T��7y$9��Fr�/:�Q�ݷԕ�{%p�RZ?אCI7�N�ex5�$�E'�Đ��r����(���-K��{�#�6����~�d�R���mt���O�O�8s;v����Is�[�o�U/w_��Y�[͎m�-��̔���0�\|��͛p���F!��,:m����f!�x}\����o��a�:�u��Ęࡹ���B+����v��N7��m���E�DZI�0�P���Τ�uc���H�G�^WFO�j�i)p�ݘhG_-?�h3�����0�n,�y��XIT�W�����y��N(� J�+��$�
G�m�?I���\u�ϥN�F�ϥX����_A�}�V�� ,ʈ4~�.g�8{�	�`���V��$��l^O�������R� �[RvK��n�R�	�%��ɂ-��n��O�׀������9*
,�xN����@�H�倅���w���7��.(}Gqa��.,�jl9a�+9|b�p�7�z��Wǐ!��P�� �������0�h~����#��^�~�F|H��|�q�|�]�Lkɗ�<�6 m�"Ӯ��ⳔBߓ�k8���s�%�p>;T�L�q"s�ƙ���o�pnp��Q�ѨWL�Q�@N_���HL�ۑH�����z���P�̠)��B)��@e�q��(�n�\�����W\�I�%kk�"�s�R<2!b)������/�ZC�+8��#P-�kZL����uR�E^�AA���d�ʾ��(��wt��ˀ��	�|#�Pe2j�,�)����asZ����d�0����#&�u<�ᄋ�Y�*��t�t3,kwGL0�zn�WbI�:<q��P��\Ў5׀���GXtE������Q�Z��#1�5��#K�3���3���){+cc;q�yd��"ov�O6�cH	����9�0���Z�Ӕ?���y�V�����3��~!�U��zL��0�<��&MlX'���
y�|qi�_Osd@�֚��C�K�KiǱt~�`�Ci��0��x�yH��������01��g8��^�#35�_�~���Y�<P�P}O+��>1�=J���0ѯ��io���f��#����?1$w�5-��BDe�Ã��ւv'~�W�)��Q�L�XH3�)\U���p0V����q4�.l;�-��l٧����;��݆Ru1��kž4�
=��6���=~����?9�V�QK�^��T�-�6��(�XaM]P�X-�=e��p*�K�49Z���	U>1�3���:����%j��ɁY2�Ļ4���O�^�g�a<��gJ���Q�^�h��l��j�Q`RY�l�1�]y��+���{۹	�m.�Oq�)�0 !�R@�@(�:��ORy<]+���1>��ݤ�j�R�ܖz��!���}�:w�*�}Ҁ:۩�m�X6K��!�#�	�7����Q3R=��ˎ����s��ٖ+_R�qa�j�f��
(U���-�n$\��b5�^ֺxІ�70��F��lb���E�y��~ (M��i�E�o�����ϚS^�J��]ȡ�I
��q�q�hc��d�UlI�@v�-)�\$m��:��K?SrK�M반V�V�A�~__"����K�5��~�eru�9ھ��g�_��+�A�'mY�/��o~��I�%�����?�G\���Κ���?�0��p�v!�Zd��`&-{Ꚗ[��������4�P�+��jF�a+��?��u!ra�Y�~��u�ǈ	嫺-Ř��mڳ�#Z�q��y�Y�����>�Y������ת=m�U��" �~�K1�*e�u9i�#6�kp*ީ�$
�F&&H��'"�t���pp��Q��-0zuZ�����A ��u�`'nD��(t���a���1'�hY�Jӈgl���/.9z(�0����m%�3�r\yu�<e��^��mlcv�������=�a[�K���W����!��|Ux��z