XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Rk1E'MK@#��^��x�rǷ�#KV��R��%�ܭ��-K�����o� �eܤ�%#Š��I���B�p�b:�)J��C����N�io`��P��0
���ः�"n�\�g�ʽÄ5e@�%�;�W�DJ.Z�ZOa�(b#��[AJ���u�s��L��k�
ŷ!��?��]�d
��µ��D:��);@���,��l�1���#/� ��E:f�-�Z�yudB��PS,�����&�#�;V�(o��m�KrK>��h��]��b��H�&\��v	�<��<�����}�F����w����F �|�U�/�7�G�A�I�*kO�`�&7$��rF�+����v��!P�oixСYGo��Q���.��.=
��y���sfY�:��P:��G��|�B�&vź�C(م��(�U�j��5���x5Q�k"b/�����ݸ���4[R�F�C��@ך_+5J(��7E�A���˚�S~K�2c����W�<�J4�>��������3�Z���_.��"����o�<�6^˓����K��?$��î)��Qb���6^L�ѝ��W�����e�=$���U>m�=$4_[7)tt4^A�qHn�z'��ջ�^$2�ī�A\xX����fUS��T�f���U�D ��Y�z���L�$o��Gcq��j%���_�^�&2�E�uk�:���螺����]4�W|S����8,�y!UH���h`��s��_d�/&]DzV��e�����ʅ�XlxVHYEB    6014    18403%�AS�E����!(��pNu�靛�Z�T������= 7����nTzv�j���P6��v0�V�Jv)���qbO^D�Y�Wʟ��b��m�~�%�Eg�������0��b���"}t,�sy	q
�)4��Ie�Q��#��;[�^�˯�H���0��@�o�y�)	��=�}�D3�&��P�^b0�$rx��C�ė�%h`b����'�l�c���p�C{jm�MB� ���2%��5���ъeK"�'����`�Q�{�jքxR�����72{�q�������>J��#F��t7�o�F�Z��,t�s;&�a���/�����f�T)K`z��%�/��,nh��9GX�P�	x�7�r�����U/c���R�
���h�[��20�@�b�i�s�ؘsu��P�T�u"�b8�߲�@xhn�TJ�:;�AP�!��� @ �gXP�c\�@0�p�m���z� ���Tx�5Ŋ,)�!7[P,��T�~�
���Zݜ�3yh^��::Q>�aI��(���qhȕ�4�:����7�U~�)]U�IF��T_�?4J��-?�y�g���
�O]�"B��<�A
�%�j�;`6/+ȴ����vvQ=\ ~*�f���c¾��r&N#�,� �p��w*��B"�꧹���Y�ex�IS�6wQl�"_
R삚�Pa%�tJ�mQ&n��j�h���6�3H��DcA�Su�Ў�E���,��S`�]�H�Pk~Zq"d�z, *�#q�����D^p��,r>>��7����N������j.�k�+��9%K���>I&����&��c�~.��3��������[쾆��]��U�!c�}B�{�6b��I�p�u���l�j�Cۍ?x1���)zR8-��5:?%��g*f�u��D��O�[0i�6X��|�X���[S:V��rb���{�vڿP��G�z����w4�����>�Q�D��5P�:#���@���p��Sr9���r�l>~H���j�(U�@�m����ք��^����'��?eZ��;�E��PA3�!-!��ys��M�l�����S?�i�( ����~�^�� ���շ�,�s
F=�1#f�na���{WLV������H��K��i��Y�`J����?{���� D����\6}��g�i�L�G��W���[�#���,3p��V:�C��\�s����T������@��t(,�i)��ɓ�k��^E7o�@aC۶��d�cO�ݤ��Ni��]q��B���In|r��� ΐ�K����	�T5�RCNkn�<��|�DwC�?ċn�G�:H<ԤT��m�o�i�S����<N�ɺZR,~�I)��*��� �P|4>x��a&-X��o
�����Y+����Hܹl�|�
��׮�Y��3H�̄��<� C�����n�4��&K���J��}��[;/w���N�������6(5Q��>�B���Ev��2�4�M�#��,�h~�� ͻ�Y����e�鬁e� �z�p��(԰�ʔ�D�忠�h<�QȬ���d���ԁ���j�"к���45�p�#q�E��j�l3v׉�c}����cN�h�<��go���j>��Y�����G�o|��RA��3U�<ܢ��+�tM��p�*�:���Ԁ��uB>��4zGPD���}M�ǋVZ��S��mO���f�.X��n�18��fqs'� � 	�/J�%�Fƥ�?-����4���j�#� "���5��N��8�O�F��1"ͭ���!:�hߣ�iT���	3�r� �"����TJmȰk���n�:١���$c�>;�l�"*?{�����e��ێ� z�NM����cޕ��(��Xu~j'��/��e̤�X�H�`(��'� >�]E*+���jaFg��x�������+oDk�o��{�ѩ�0~���N�E�5�b�+�?)����t�ny�����.�����g͡Ṁ��z~t(M��i��;β&j���k Ʒ��k(Q9?���9];�ʹ����\��H{Rﳖ�����|cA^�kD�WLU�L,��P�"�)����=����f�q��1�ū�]>8�XMq>"I� �B4U�NN2��,V
���S����ʼ�%�fFj��5%������:��}|����w��Xf�|M�6-�	9�F-���3ٞ�c��{�ﵵ���������P
^W��[S��ƚ���h���g������~���_��%��V���85׋�ĝb˥�MN�2p���q�x�}�`3��K!�#�F{��o{K����J@2��P���(���b����]뚊�J(����ۂ}r��1ǳ ��-ܟ0o��w�1(g���D� Ɏ��a_�k�u<h���|����Q��;�W���6
�.0�pN����E�xƹ����c�Qx�B�p�Qi+��1m��eBIdFpf��A:��ɂ���6;��`u+���w!�-N98�QK�W=�7kP"D���)'fS���:�������&<��|6��E�z�(�`��\��zX,׵z���A�Nb��x��W��QO≄�����"�1�FK����i���	�N�l*PgЊ����a\Fװ���?��+BN$�x,���C��鍕��]w^�	�4�Ǽ-j�o2U�+��c��K.p��U�+�:2��Ĩb�z݅À�.˶�-}��h����Xn$�+���p	q1���9|~n���R[/�$�愢' �;�i9�k��1b��c+�B�V����r&���A�i��g��ǘFz$Z��BǏsi���Ꙭ�	y�����r��`"�`�H��/�xq:��c[��sT9���s�c�y�a_�e
:�K�piaa�h��=�5i�Y�I��;�8"l� �1ϼ����aEL��i�s(��M��Cdnhh00M�H*�E:��=۵��s֡�0��>����
e��g�^����r{����n�����Rw,��5�N�a\w���	U�|�%�oo�
��oC1�c�8�/����� ���%�)ŕ2U���x	��0^����7�O��ސ��H�V��*έ��<x���F"E
�Qq���y��������
R�.l�y������>S7n���	� �OmT-�[Y�XQ��a�66h���,v����Ӹ�k���YZ�+K��{�1�cu�(��{H��)�h�����"h;٨���j������G��� 
���ƛ�=�V����,��3x�"oq|�}E��C�~�T�֘]�Ј��]Le%m���*�����a}zǒ��������� 1`��ݟ}�����������R4�y~~g��g���ؚ�؞��=�l�4 �
�x+��H�0M��w��quʒxg)O�Z�w��4Y^��Y�X���}Sm�"YTt�E��}q]\����^e\�^t	�i�(���������D�R���W��􏩌P���@;u~�+�ߺ`3���qm��� E@=N����������\?VgR��gZ.r�"�9s'�K�1G|���!N���_6ՏZ_͟<'h�aI%l��d�,\�k*՜�Xu��~nnA��G:���@;� ��<�	sW� �-;��V�f��RaV��+� �<Ho���^<@w�� �Y�N�6��M����8P�q��b�T����?22A}�����n�i�i���ՙz���! ���?�7�bGU�M����q"�ڟ
 �3F5 --�Ѕ�RM���Q͎$lO]�E�{�%*6�F��l)�����w��2���c��6�^�*	��T��V)$�ɟF��'P���8'�QoD-#^���y�LL*d�W|0@EB����L�Oҭ����?k>�?P� �|$/�W���f@��L/'K8<�!R�+��u��mT�NG$��6�9D�+w�|I�U�\ޓ�9mA�H�ݓ� u꿽����0�:��*°W1	�h��t,$Ѧm&�h�	�3tCV鐲؂D��� '�NS�>�m�2��b����R63�Q����2A��.9Q{(���"Z�xa R�d�yK�V�����[��"��8(��G��[�0�CX����x��s��o���S�R۪ؖ!SZ9J]m�jH�)�UN��I0$�qȭF"S�ͩ������I�6���F�v�4Ag�)+�?��kS%'�ۻ־翀F�A�޳��jo�4����ϻ��8mN�j�$��5P	�̍z���"�V1X;ѯ�
��ݯp�2��s��&�W��c��P�k���m��-�5��%��\	�n�^��{^�&��ݵ��K�4�^��17� �������K6��t)W�0�=�e�� .M�Uq��ar}������j�Pa(�@��*U���T��=5�-�W�	��U�V��]U:ֆZ�PV��[w���TAt`��i�t0t��s�ˋ�dFu�n�,��%7 ��6�/��s��喻ڍ�	2���Іj	��b�A�p�w��"�Ss��VW���!��S��hֹ�y�{�N�����J���!"�D��
�����' ��]5�N7�^e�)�>�����tx�3�+�D��?�(�I.K%ю۰
�P6@ޚf�$n`&���:'g�Ƚ��X�����Tf\�;�F��Q�:��� ;�"�c=�{��C�^Cj�һ�&?�1��@��Go��[k����_�\�(H8�w�m��6.�zV�s�kF&���i 3�^?SawS��]��g�y���\7Ȉ|Q�p��c�"O^������d vΙ^$�Ҏj�]p|
����$�驗�Z�I��x��򪹳J��HaIq����bs p�%!X����*�|�'�>�m�O�����[c�ϕ�o�����O��pH���\+<���ͳP+bڶ.-J��^��K}���5��y��|��-/,
�7a��î���qo�!�Ok>�2	1�p��'�rP�5m{�ݺR�6,V�͓2%~�5��݈ǽ�q�]6�Y>8�]�%��a��|�p3/RSHG�c܌����	����풽a�xfXcsC�#><��od>J􆏨��{/@?�e��Q����zPUө�)ӹST?�
�	h.��E�+$�Th�K��Y����ݐ��|P,�*���$3T5�=F��jE��؜��G���`~u2#�=�=Wݞ�ㇷ��l(tWca�w���9|��,X�B���62��jVp@�Dm��׆��Ä�E��)Q6/N�Z�c�<��p�&����(�����>G�{�&�0���vg0L�j�m�K�<S!5�B6��/�@�����N'�� �Bn��>��]c.�����e�2���g伍���$D[gW~/�	�gF�$�դT��_��c�Q������
����^ߢ��,]����Y�wY/�W{A�:v#��%1w�ƶ�IЋ���W;
:�㪹�[�wR�H��)E_��CzÏ�?]d\&@�P�'D�8�Ϻl��a��ҕ�`�~~ �@l�Von�>H�N-�|C}�Z:;���c��k�C�^L���J���}��G?�]K��D(��w��n��?�Y�Eb4Y� �������t�dr���Y,gӽ��>��"���u��,��ݮ�X�SWr�8Ȅ�&K��@ä������C�:3\?���d�\%��.��*!�����6�mK�՛�B��I��K}g
��5q.�D��l=��A��
e��ʫ�P�$� 9��M�H��-�'LPU'���(���̸�.黾]�Cr�����ru��X^ʽ�����wx`\V{0���+#7�S�qN�M�xӜ�)��P����ImT�"B�ImQ�Ғ��B�X��(Ƚ�uͰ����έ)/5"C��g�o��-1��oU:�u{G���
�̎�<G�K�~U��C����
o
K�F@�(�䐌�S6�B���
�C����F/����4��Ȍ��c0��_�������EF!�<4l���v�t������o&�^�$�R�C=^t�8u��N�k�Y��T	����` �'h"x��s��W�ee���o�J���`(U;��g��<a)����m���:7�9�,Ɂ�B��\�B�l�,��=�0!�E��;�͝��Ǭ��67