XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'����=�ҥ���[8&��^�T�W���P��B?%��i��d{eD�'n=*!�t����y�MrM���H� �YSK�{,9���o&��e�~��׷��mU�D�� �����j(ө�	�>\>*v�A����7��I�N��̦��x��7ip�44e)��(�4N[\h�e�@^R�:�<���-P�.��^ ���#6�����G��z�,�#��!�l�������Ύ�mO� �b��a�X1�Kݐ$�|�����xiA-���@��
�)`
U5,h��(F��}a8^O0UGK�$'���-�v�8���>��Gk
;3n,�_�J�h ���𦾖�k����L:�������9k���6�*�  ��O�"�9G�]��~؉���N�w��୫���5���hm�|$U>ǯo���.3X6��ql�ۦ�Ԃ�90l%
��Yn2oG���L풧y��0E<T"Ms��z���|ԗ��l����҈֪x9��A/�W��'YW�ϯS�$X� �a+�����ʢz*y�D�Jǝ���I@�~���B����C�~_R3�)�o��9�x� �DD�oV��2�S�Xp	ˌ��-�W��A��t��R..�Uе�5��0�m-y��}�5��X @(!��2=�a�J��ԅ����vׂ�|�t�B�D�٘:��T*7���(�x�Xڕ�n�>�y;����[*�5��ŧk�.䄀�=��Sc�I*�<�ٳ�/��lPNXl誨9�Ag���XlxVHYEB    a037    1fe0���^Żǃ�bJ�wY�N�㶐"aS��n��� �_��XR�>s����c��,����Q�Ц�WY9á~bt��������$�(a��3k�G��V�1��T �#�����]�/t�$ئ+0�  �?���YK���Oe�`*ޠ-?����~Bw�� B}�S�X��7z\Hy|uGf�>�-%g썡���0��_O@��\��5p���l}�!�i+G~}Ң����؍�>�m�����
-��uؤ�,r׏�~a�3'Ma@��Qk~*�ו�Նp& ��>_w���Z���5�MC��%!��c$�.	Y�	�<�ʛ���7մ��@0���� �t�*ǁR�t��h�غԡ]�y>P�F��W�(c�q�QENll�b��[J=�8Js�UΌ�Vٹ�Ba�"� <�7E�~��؍e��^gVPK`EVURnb�f����?�f��w~�Y���]�%1���:V��O	�ɶ������/�m�"���^ei���r���D�����},1��&��*'���v�%$]P+�9sv'���X}��d�����K.��Ѭ6G��
%!��/MYgF�r��)�5cݘi���%vn;���A�$Z�l�I�=ve4�̶<M}u[`%Bn�e )A_�����Tn����3���O�m�zå�߶Ӆج�$��@�KJv����)��6����|V��Hn.P��3y��r�p��	�o��&����cl3�$ԁ��������?��&�
����bKX��l�-i���Y�6pY2;�)U^"��Ԯ�-}LCU��c`:�D���$���M*��q���TK�6Ѧ΅ӰC�}�1�	���e�Q�7��L6�pha��|jgTI#�HЙH�PvX���;�/�7�)��J��&3G˥��ZY䔟��<�f�v�#���m����y
{�Ǡ��`<m����, �g�腬r����"{2P�����%$V�g6/z�.0�*����o�X����ZGg䥦��$y�B�&�}/#�)�G!ǎQ�ÉL�:Fv��)���r�`�P�I"����4��<�4�b�ƒ���@���'MuG;���dB`����.DoZN`63��Q�����wH���F4x�B��}�O�ݯ[O!O3�h�w�&TUۙH�?{�g�O}��S�2�/�h� �P���1�I#��U�D���n{����A�ϒQ ;<�O�ڠ��@��,�{�����n�/~������!����x���%�w@4� @$`s��O3U���R�_�(E@��7��$�v��Ԝǡ���X�!,W���Dd���M�ժ�$3�]�M�'`�SZ��d���\t!x�~M7����a1;~Q��24V�E͋Z�
}9�����X[��|)�E�=;������/�/Ĺ/m�'���LN$��v5�3�����p�}h-_��♌��P��t]���gH��`��lT��d��_��.8&�� ���"�a-�<
�b���r�2	9�j�N���/����0��~�v�8�ޟ�#󂢦�!ɱ�kGe�����4(��q�:�up��a4Ks�"�J��FJ�Ø���h��O�5���c鶸������9y�m�<W�����Dܒ[���[���r9ll��ۭvj���Δ�8���,��'�~���b:bj_Vxa+�4m�y�IZ�$�%5r4QG������$��Ҧ��/��>�Kz:�;�upBʝ��ޏK@�j��{:�*��rq+>��o��`���M�3��������K�Cr�P��&�o�� �j;��^����h�݉I�H����xW�%4�x�{Q�9�i�.�F���S���������`���0�Q��ߣ��Xhs[Jy��Z��2|X��-���,\Kԏr�hh�A瘱�>֎����(g��WEuA�VaH�9�Y6�AXcs��?I�Ԣ��1��cj�Jg�x�E�k��쐙��?5v����5����gET�)���Pg��\n8P�q�ݦ�(�;F��7��I}��P:V��K���鏎�3�1�<\c~Cl�.��|���8Q��ma&W��K�<}��lv�[��>�h��G�	r�����*�!�EN}%u��#�kÓ�E��BY�%r}�3��Z�K-��O� �s�<�"���*D��U��L�#7t2�[��ڥ��$k�`���>�<moP��e �j��Ub��J�[������Z���ޕ�$tR�w�i���@�'�X����r�893�i��Ý̠���H��X�o��U��BՏj[����V<�Kg*�L�𯔙q�=A���0��A�h	�,�8T������f�����)g.� �@1�y �l�'Ѩ��SѮ�Ҍ�b&��D���	M��
.�+��$ϴ�ACf�A�O�y�<���xJ�3^Z����,W��cMj � �?���Zo����*�P��0��5:L��i0T@��nB�Hi�p��
�lɪ���-V���]U����,���=;z��Y�u(�C�N���Y�������廀;t-w\�T���z�-��qZ
���GH߁+��J�^̪�=j@�%���N���Ӆ�����hբo��R�2�Fl�����nJ]�Zϵ`.��,�] <'J��Z�F@�2;�M�\CW����Q��ZZ*�%Lf�2&��� ��*��*�Q9�V�"u���q ��e�W`G�d4ob�����"����&�B�C�A���w_�������hf�$���Y�'b>��r�G'����0�р<�YN�"~=<��qЍ#kTs(�8̠��m��X��_MB���ܞ��	I�8�� #]�p��4`n5*I�V/\"8?H�{d�@���[���&�K@�$j�����|�sb�L�0~���en�H$N�*��|��P['��0nv��5�����ڶ���q���9��D�����"1͝i^
rJ����u�+N�Vڴ	Sr>�/�>q�1+��C�̈́g"����z�g�0 ��cB��U�<��c��=��Վ���YZE���@6�m=4��*wUz>�g}��Z��]��$�r60K�V{��K�W��M��d�>;��A�yj�5<��8�X�_\�^�X� �����uĔ!��)O��ԃ���,L�l>w��)'�a�-�e=�S�u�=$��2s���g����p��T��rO�ca�MlG/�2��#I��Ii��ScWT�'���!NX�t��?@��c����wZ/i�Jv6 ]c��C
�|��9�)�nC��9�S�Ⱥ�W����X��5D�	��K��X�G�ٻlW���f�g��.d#Ɇ���Ejw3�h����3#`���J��M��p{gd_��M��t�ڲG>��.��2���]I�?��ި�׫�a�8���)��d4Vʷ=���
^�\��]���M����
U6S���'_8+v�	^0����M�b�n����ޝ���a��ު��Z�Yڣj�S��U#KU0���E��"~]��7.]���W~���@^��ʹ^���)Z�/�1D;��r!�d"��h�����q�P�J��i�:��ŧ]��Ҿ�F��`�=8�֪��J��=��=#=�Z�˩�W<h�l��u�N�&W��5�2�:�h�k�Yٴ��H�N�aG? Q2v[��.��N8Y`t�(�"����d�b=P�ݿ�dp�����է�q���JI�{�.�0-�ӕo���wɵQ(��`��Q�;�=	�|@��J�k�D�o4��0ʚ` t]~�W7����$ԋ��'�̘���/k�':i�'��@�\���R^q�m$����I��J� =�f0���	Bv���X�5�iLUO��p˅ع��;gdc���$c�
��ט�$ZL�l| �؃{��]E�5vD�W�����?�{*��-#�,ꦫ�5��j(A���W��Ӱ\��W��N\́���p�ͫ��>E�
D!N�1��ɩ��$_�e�������3���=���}t��b��R���L��'��kcA��a���5���d��1�7����%_n�����2�&�t�6�����C��;��V u5L�P��/P@8���g�S���U����+x�zs+ޮ[��;�-K�s�!��
N�np����2:�.܅��<!5��4����.S����^$��ߓ�?,:uJ������=�GU���'B�ç��"y5��i�'H+�*�B
�G��jv2��g�A�M v�S���[	���R/���W`+k���#_�Yn�r��(�b�?�<��^�8���d���h�?���of	�;�o%yWtj�.�z��F��8��.F��j��{%��#�H�.�Q�-�<�ҝ+Kvag��p�u��x�CÒ�v�AA��@�J�B���������˼��<��E���w����f،�Y�zYN��d;�.#S�MW�=p���53�r�+��[����s��]͸�p���`�!s����v�s��TX4�qk��;�)�='�񃷡�nn��!@}��b)��2SNso�c��C�8ݜتU��b`�-3n��9�
(bQ`��jܒ�u-W�ѪK��=��v.����v��2Ω%5q��6�.��7�9�͠w�ns<[�]��|�F�%S��Ve�����8��9�僾�0�ٖDT�q�s���x�Z{�_s8bZ�q��\�5�����l�D���g��-�	H�I�6SH x��ΎR.�'mW�b����@w�o�oB2�!������{���vYa���\����D�5�E���4lk�ė[�{4��P�MJ����L���b��\�4e�t|&m�z/��}�ơ�n,�8!,j��+�o��1?�4� � f�z�}	��	��ݦ�����ycr���J�����>7���%�J=��,�B�"��b�+�S��E��juV@qVV��>�O��#����9��2 ��� pוC0
�����>/w��sk�n�>�@1�� �Lj%�|����g6+��Y6�b�� �?��v�S���Y+52�S���x5�~��)�����K{Qs<�O���P��J�%�D��mz��4�M�,��!�4�E�gA�8Wۖ���]��`�Y������l�N@L��ͻ���������$X�ce��T��Ѝ��ʸQ�3��/B'WB�G�$t%��Ŧ9�d�J����-ba��i2�Hq 켥[�`���=/0��W�M��
=?�)0�ʔD�/p�e����9�����i�o9 ?��b=��mj��a �Rf����	{�1�Fuww'rJ�%���<E�4��h?���3�k�6�;��j0�R'��0ju�ޠfE\s�B���D����2�p��aN�[]�U7�9Ŧ���#e�xu�-�JYQ����[�,S[�(� 	C)MMլ��#�8��������?�x����4��֓�p�S�}�bf2�|�&�-�q����ű;��6��6`އ�͇����E/�)�Ir��?^h"t|�+]���8��L��N���o@����w�����)8#u�TW�d�8)�8+�s�C~G��Ɯ�ݝ�A���C��A������z��0�C��2�}�S��ӳM	��g�V՛J�9�'��!>��!,��u+Z4�I��!5�MلCy� A��A���}<����q툎Pw_/+B&�~��j
_�U�Yb�U��5f�r�%�a$M��a��aW[qD��&�!�V��}�iR�Աy(�Ae8��&i����;3&W�(Y���Oz�Pd$l���N d���Q�\
BB,E����"����:�x��'�$�C��EIB#��_��rStm~9��1�J}c}���N�AZw8�\��/� Z�=�(��ރ�
�t�kXĭ�\���IѢ��v;&nኰۋ��G���`�����Jl0��@?^�m���ћ��p����͋����&�<ۧA�I�O�őTL���s�ߖ`5c�`ݛ|E`���*�ЛA��;{�1���1�s�ӷ�0`����kz��Dѵ�z� 3�v`)o�B��7��oq=ˮi���u6�6��v��Sr�D�G������fi�,�� �?��µd|t�olu�Q�\��a������~s�����V��93A�|y��M�|O��}��;w>f�: �v�wV�q �>�29)g*��� $����6��4c����W��:P$���o�uCb��7l�bK%��r��|��	���=�G��٣#�~��Ѹޙy_QqG�x���y��A��'�b3��Z��_4�h��j��
B,2�tW�+ؘo���g���������T*���Lg-���l�
��n1�Tq�8�b�,:q%1� �b�f�wRAW����x3�x�&p��e�`�����x�)9���$cfk��$2u�Sַ���e��[���ΏJ�+*����ُ]6���$#��+�H]�B$IDC]|�MxD.��Z��=z�*�(�EȂ�-ZG��U���no�&5�K��J��|D�e���];��-c���� � J����Y�-0S����'A䤇�-�x� 3[fe׷>
&�,7�U@J�w���ќ�@~�-�L'���A0�A�i��D����"��4p�p�d�'LN�
�(��d@1�j48(�e�Oc����N�9�7Nm�S��s��ݪ2��O�es.ԣ2��p �A���zlN��C5�Qe3d�+�=`�yl���o��H�v;p��J�Te��f�\"H���w6���Ra�l��KZ�`��t^l�Y�<F$�`k�q�	�g�DP"���@��f�ڶ��7�&���5δX��`}�n�@w�
>3�������C���h�`�q���Tp��	���!�φ�"�C�<AM�;���h�	rB��@rc��s���x*+��T��94�7�#�L)!�Ʉ.g������������0rx�����3�~0�X¾u>�i�F�7("�����m,E��=t�0��=��#�s]sQ�UAt�fZ�v��;�f/@$o����6��.b��|�A�'�6#G��q2����{�}��.p�\���R
�n�<[>�qH]`�W��G��fw̿{a��՞��R����f!'�AH�O�q��p�_���/s��� W���d��?�\o�q�='1�<�a��%h�F�XS�ob�7��ݻ�Hg���/�R� JĦ��V�0����X�fYF9!^��Np��8�e�۸�W����h,	e�	y7�0Q�8���.���'�$1(/�l_�+X��o�R�X�[J��Z�A�q��-/�>)+p���G(��X�f�Upc
��Z�S�9�\m��!��\�U�w���;����	w���Z��P$��&`������XXL�!ɸ�R���Zςܩy*�_:��Y���6�V+�>�� b!T|�R�s%���#��J�϶d�{���#fp1�z�J���oȗ9�-�ܷ��~q���R����� :����]3��pt$/ӫ���CI!�[��G�[b�8 s��h|4Vo�ʡ��E�20�Neh��{�a��kF �"�г����.�(�Oi$�^ ��Kb�	.��U�|��v�<��l	��2fa��*��R�_ȷn�������򨑩J�Sf�tv�w�?����T�o�ʧb
�O����?���È�}A<������+�"�����S��ޢ����GgK�ޝ��Dz��= ��U�E��J6KmՅr���� �ؔ��7�:�Lt�y�T��I��Z�l6J�����n�yy��{�Q��#���*�4Ɂ&P������f�I*f�59���_�tz�N�;yOl���@�ḿ�
5x�f��w�)]���o����;��C��ID��Y�:
ͧ��*�H.�`�w�]�2S�a�^�1g���WdW�2G��:M��op�&�	kM(�Vnn	)�;uߩ�=��;�ޤÄ;�fS[��*��B]��m���<���$�U������,�=�h�d���({��5�UQ��s�5rL�	
[h