XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���g�i�z8Q1(v���4�%��;?���2��NZKK�)�h ï�Ԭ�`�U�&�uH�!����y2H�h���:`R��q��	Rܳ�$��2��p�fֈ]�cE%AA
�3�|���;ۜ}~^-�j����N��B�m�/`ɓLF�]ƅN?i���(�RcGFn��Ơ��˟�s@o��:F$|��zFؘ7��Q�K�.�Z��P\�\�� K���z��ҝ���%auu��"��^��m�1�Q,�Oު��F��0���D���y8��N�ݧh�Wa�w+-#�Ө�
��F���*��n|l�[�G�<-	�OX�i�dLU���0�m4V������k2�Uܵ�R9\gL�!���u��f�̀ز?P��Ê
�h�e��B���m�E	�ǟ����]~3ű�VRf5�:_>�Q�i��z}��.��D�R;�X�Z۹���!���������~rܾ^�y���{Ęv��Q�|3 ��=��B<���ޣ�ۼN�:�^��JiK�0�`�'�nd�:�>���9s��=���V���o7`]����WDΧBO��|��@������U���[����T��z�l�x6!4�܁)��ͯɒk�-�?�C�c�I��؉3�,c��*�g��d�;�x|HV�-�T�,���H �e\��FNQ�$�F�����!�����z�+<�iǭI<�rnE:F��yd� .�Ym��w_,���-��t��g�Hm��s_��XlxVHYEB    95d3    18d0�1"�U��$�-J��^K�j_���xz�^�8�,�Wȥ��Q���X�A�Q�dRb��Xr���U��m��}�>};�KVhnA�3�]q`@��2�Y���t%S`��DQ�ֈڱ�	& LFr�@D�.8���HίiAB�H�]+$k���y3������F�?���������ot'��2l��|�+}����u��!nYFS�yyT�s2���l��Q�0�w�:|5��@�x�gg��N4��Ѐ�`��KjSW*�a�h݆���\�n�z[�t7�e���MG*�T)[�:���:�߆i���`UAZ���ٖ�>���=߭���7F��%Y�&(C�cct�G������/`�CL���Z6o���dH���߾�(u�؟9 �'76�������jN8���>	9���S��W�S���/,�uL/n�[�@���liMXBX�-䦯���.��z:ihdjW�q��+���)����<G7�κ���C6�5;.�YU�}*C�a2y�2��B#	���(X�"!� �����*�:�e���O�3�����f���F��-ء�46��� ��R���WE��7�j��>������<L�Ka���90h;D{w+��Y�L�A���.�oƋmC�D�x��| bSkL-�pkn1�L�g51�]�#ҳ�.mX�8����n�`�� Z�9�\�睽1��DïB+h���-�.��0���=)��2=���(G��F��*Rx��@V��YN�q��uӖ:_�Kٖ�c�~2��)ZEU�r�Xm�>l���/���G���Nqi���3](��c�<b]�P�9�B�|���2��$����@�q�f�Nt���_<�����y�͙��$��Þn�������Fm�6U.s��e���4s<���S���u` I:'�9y@���� f)e���D˘*e� ה�f�mtj~e'fj��r����I�.@�~p�g�/:��w� l���[�0��uG�Tt6�8n���eJ��|�\U)�����CAj�#,ª�`#��	Ē=5T��^�-�O�%׷`�ū&��;��a�*$��^���
.A�?|��0�o�S�����Ɣ�o0�ԏ"�%��<�kv4�r��eO|�+@��\ÏG�n��� �@�t����o$p�i����=�0�t����B<�Ģ�e��	��ܗ'Oo�jMP��jEɐd�K)��EX��d�LZ �D5A6����/�m����u�h��q*�Q�����d��Q&�f��W�O�y����r�)w��`���-=������6�8d]�����Nh��o{��")w�q����Zqj������J9d�+4y�~����)�"�T�n������G��K�8��X�T	��O��6����V��Nu��b�d�)ZX}��<0ݒ/ !	q�gQGf���<%�E�/�-���V�!�1߻xAΉfJian�ÿW�ef�I�N�p�&p���vgh�VASx R���uG��Ԇˠ��R��S!�Dj��/�s����C�ٲv�HLq����V�����#��wq�+<�3L��?�m<��O	����f�u�LN�#��^���O�Ӫq~�i��巶�m�!�{��"��N���+�Ϭ{I��[JnV�l��Y�\[��'-2��M0�
�6=���#C��J�?�clz�<��5����:���v�9�!2�
��ۙ7�L5���T�14�����j��HⳞk�r�$�w�C�$�Me+�߃|~�y�xY��-W2CgY^�^� 6	 K\O��$�)r�N����B�e�t%��V�|~>��[�(�h��o /����"����Ahb�``��Ii�a���w���%�<c���B	w?�2U�N��-�NK\@G&��8��A�W +vd������%S��$�_\��I�g(�3�(��P�昺����(:((D��j(��aM�s��h̕��G8�v��y����&�_�{ �/����g�+�G���5c�����4re�򇙰-l�%_���l�2=y� ���Md��Ǻ�#$�[� a�����5���:܉�񆮋�9�%���	W��Qم�Z	oe�?ϛ�����ɶ:y���KM��`�ЗM����m� ��vJ�������Ju#TXb7��3�[�m�a���ך���U�HT�čg:l�ƣ�7���6��^����l>/����ޯf��(=�4ϻ�̓�Ue�V�σ���I���uEN[�uWTj�ܜ����u!����^4_+*�;���8k�)B���gf/wS��$���a_p���F���N��Iv��L�EubF����>91A0Heg����:#��>�u;�ݙ@&���b�řz�
�m������Hա�)}�p\hδ�TU�j������a2�g�sEol@w�j}w�4��jٽ}-�'&48�?�m��_X���=$u�,@g�|�`
��^�l="�z��"6I�L3���޿��d���Lʞb%������ �HJ��B�V��,��'��ǨvEf��.Vb��#t�:U��)�,�q�ա�?Zh��Ѱ
&���,f3�R����v5�i��#�_L�瓑��`�ԁ���l��S'�����w��ir��_��Xsfh���P��Ұ���H����<n0R:��R3�݉�|�[��⢊���G�C�h���WYN]�oyPD�dcb/��
��(s�۰�!$������d�� �o}�-��18;6��Ik�Ns�I(�-	"�,�i�P��y�Y����z��r�n��Ԍ�c���ݰ:0���}���x�ڭ?�ж$_�Zs��� �~����P�fa���*(�/�g%��o�������C�IgugX,�8�ูp�4�r�w%��µ|����/w�}�H��mM����?ʊM䪃�[��K.
�@`a!f�͔aT!��
��-�*�Z�`�@�(ʜ�$��X�_����9�T�~!����26�zm��pf%VZ�T�Y�8��_2>��~��g�,WxAD'o�:�fr)��v�x=IQԻ�
A�A�OtR���F.�m���*o����C��BN�O2ɯ�D�l�ŁR!A�d�@P���:+2�N��^�f���| 7��$�Y3����\�I�i�X'0�K5�������jխ0���k]T�@<Q��7�����������{4���O�<�������L���A5,��Ѩ4���e�Y)�}���������M�;I�P�O�b��u'�f�cU|�I��Ǟ�gy���:�Qo�S�6�_FQG��M���M�}sp���@=s~����J�D� �e�(���J���
r��Dp�*�����d�tn��A�F�(��QbD����ÿ�z�k�$q�h�'d�~"� �ס�۷	DJq�[���O�R71���|��dx~�X��7�rjd4ܝK:��`2V�ڝy��n��ގ�wb��<ȏy2��'U�9�������ď�M�P�]!Tc=�����3aC�TKvT�r�,?����;	dT��rn���"^�NT�0�:6o`�SZ���aZt8������� �ɲ9�r �V���!98#�5n���6�zȤW���Fp[��̰0׉C�WK��)��EY BН'Sg7@=�~�������G��-AD�cV��Of}�s�J.
��]RR3�g���m�T�gA��K��ه�`�����M�/4��F� sgXؘ>C�g��>A�C���U?���Nq���hȝJD�����9��c�k�(��5�]iy�`���qu������I���$F�N-!�x(�`�Ʒj(�{�e�w���e�a)e����}���9/�	��9;����-U��a0O���������	�I7�L~-����
ȗի�I-�rz^6lǄ�Sd�'��n
7�U�����",;'ASX�`�q��b"zׄ��l���Y�ީy�I<��:�{�����.��{�أٳ�)̶��'����_�,j�X��qv��a��`��ښ=�;��kW(��!Ѓ��<!��S��H!�»���䒒��l��Q�I�,���Bd���z��B9�2O{�*�Uq�: ���u�Z��)�q��hu���A?�S�Q���3��ᔀ-T�y���G*�G�<&���W����t��e�!�ې�Wu�(�3�sY��O) �C#����������y\�/ʔ�04?��^��S�����1�^����'gd��jJ�w$��F���j��kjx"�pʮq��O�"�ՔRi�?�G�Z���JT��Ś�Y߬�iD�ы� h��Q���[M�3�#����T������rR��>3-kMMo��:BV�֣�)�Yo8IJT��7��c�"����N_%�G�x?�l�� ��h��9A$8M��̢I*֛�+��Q1jF6/롮�|K�֦��Q[� ɑ|Z���@�S�4IYm��MH�D�_���٠f��S�L�c�}���j*�
�}��܎cgi��S���Z�*W�@H�ސ}�x��H�V�DE
n�MPPd;�����.�x_l�B�֛�.y�lB��؈�X�2I���J>�C���-���yjG�y�HKMf�O"i
2����ӓ?>V
�XQ1C	7�>+��q�ju)a\JS�>N�s:;���R�hD����:bQrԳ*��ר�>dLmX�oZ��{�.�^̻�o��������?#��SJx�����j���Y8v��o F?���B�
�Tol��⻡�M٦�r�	3g�����N��,0����'�-�hM�^�����u΃(vK�n:��R�L}��BwX��*aC�)��.���x���#2��_����=�O)��6�����J[7sD�RGb�����<d��ڰ�)_�����
NfZ4�>�94�Yw_I�2�������ą%}1�m�&��x|�  gPEc�Qy�l�L����6jW��W�S�U��U�[��N!�G�s�w<�x8��P{����� �����j��"ܣچ�`�a;	�����%����|HY�L)�V�U���B-->}��]�2~xq�����:����.HD)�
��k��j��Z�X<<6_~��g�mj�,�o(p|��l6�'Č0y(a;��sv.���¿Rb\����x�d�dm�m�k�6���H�&(%�?��ݒm��Qw��]+k�ѳ�<���v�W�L�B���.��
�$�<�)vF����"�tw�T��Js;��W������w��{	�n?��5��ċ-�>�xe�#�J�Z?�����Ș=�-���9DV�T+%�Z�aGQ"���Y*F��y�%(�!�r��G^x�!���BE��,A�]�!RmH�@<���*o�`J.�6� EYn�r��V�	7]�WJ�R|l����j���4���p�zW�A�a���64z�Y���lqKR�O�c'�hE�N'I\����xù�KO�QP�ǧ���"Q>#�_ќ�rH�e�2E�6�n�@� 	�:�j����*({P���Z<�+ $�ı&�E�c�{8��Ưw]�Pؗ�a�^�%Hx�0f��Zj����'�R������Z%�Smk�Zv���f(�C���5�C�b�&檴��4��\��x
IH�`��"�eڧn��x�P�ɺ�^�$m�S3�s�x�3���$��;��5��p!P(H�-����jR�m�K��ؠ������$167���n��{ӗaV�>o��;��mYKag�7��7
��*��z8s���i�}��,A�D�pGO�-�JTc)S���<�&3u���{�,�ZB��������U�-�	�
Ъ�sɑOSf�m�O3_ڴ��	.喙͚l�j���w��pZ�&td�@F�"O�睏���e[\.o��f�ɶ�ۗҦ�0��OO�)둣�Y;R=���8��t��ixs����c��LT�2U+�����[��|"z08�w��|b� %h�e��Z��}WP&���n4)��ݮ��:�3�|���� ui��G!z7�cX	��lYDj�ϻ:�$�������˃%�nܸVD����N�Ԧy3=p�HҢ�'�`�]�γXB���`HwH��������=#��� aak�m�b�����?,w�����q�n��0Eųe��^�-P�2u#��d���P�S�����No
^/��