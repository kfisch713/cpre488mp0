XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��*��,�&�=Q�4��О������������E�|��R�&�s�ЖU�p)�rP��0�E ����[2���[,�#G��*b�rf���,SY� }P�r�ռ����q�X�90��^����L�m�ǵ�dɩN��HPq�	�]&�7��ο��6nb6U����{�$Sŧ�^9������6
5��`�ݘ/�OT�9�U��K�"��_&X4V��1�m]��@;�2� 8��Ԣ����s8�ۑ���,�P�������'�N��&QPik��Zx���Q��{�iSR@���&C�����f|c.�WIi6���츤26<P)�S�Ϗb˙�࿫���|$F&ك�+��֞grGCk)T�quX���g,��u��P���'����Q���8�t�������R1����a'�E��ʿ.#�-e�����^����w����nk�q</���֍��,�UF�4��m_=�DE��ǋ�~K�c<3�b��饥�3&��[�˵QjGؗ^��r�RLBr$<�o�,s7����`"���Y�nXĦ�ׂ$��A��$2��m%���A,���L%��_�5���T^X����m��{�+i/�s�Uz���ݷ0���k���>�]�#F7��&��rj�p^U�' �F�y���;�����ۗ��{�t�:�5޲UOU���שׂ{�.X�� W��0�!�.�&��z��Q�2�{d�?�6O�;���{ox�eHP���C�gt�|�j��j�o��ɾȌ� XlxVHYEB     f6d     6f0��S��e��m݌��RJ�������l~�~�����ޒ	�� '���j��z��얙}�	R����0n�8��[����eQݯ���pN�Fdt�</���4ŏ�g����FX�2qiO�з<��jx\��i>.S���q��k�%�0 ��Q?����gy�����h���T��o�v���透���
4�]z:��KU�s䷼�>A����r��M QP�t���8[��9�˱]T��ce|�u�ys��%q�֮r��L�@D�u	TE�t�i#y�~e袅~��vO��\zJ��,�t���L�	��R�[ �V�!%2����?��oo"��C�o��@�L�.l�4�$9����iG���/�.â�T���lQJ�
����ƊR���)<�����EU�c里��"�A ���X�\^�L�o��]�8-`]#S�+�w�YqO�J� '��)�S�B+F�g A$`J�!+��'�ċnzsXI����X�	�6`r)�B�0#�Q��c@[#۽wlk/�NLn^pnU^hu����ȋrzb	����Ǜ�#s��4�]��ᩯ(^m�EW
*,Xwɡ�@6�%?Z�eJ�s.�:�
u%���^:��X����k�C�]�/�����E����85;l�K�˄���pUl#��8D��p�9��5���)���;�:ܧ��	f�����_�����M�O���h�h؉���]�k�!hoS�w7.��f�t

���'��Gj}u��9�|1W�d��1NuAv8I>t�^����:Q�Z��X�"ؿI�a4}�|;M�|�T����IpP�scK�m����q�1	j��_~���*����R�b�p��jP�K˷V���j�SO��G�E	�t�ߠb��~���h���u�+��A�6�~�l�bɪ(E��f���0{l[��n޲˞��$�;.���c� �4V(;�G.�/�뼵h����z�7�c�;g�����L3Ֆ&F��0��K�^*K��oT�Hyl��������U��*zx.��*����l�5�hD�'rVr�m�؆i�5b���S��1G��Є�5$��D\m3�:��{�x��.��3���q�95姲�s%�Cmn�W�AD�z[uFY��Ь��������n��	���K~�)�s8l0���1��^�̈́�)hz�HB���Lv���GYfu(��J���S""�S72 ���"��I����\���g�n|�f�~�T�F�[�lވ����+�o*���� ��b�����ϟ�. #�Ӧ^�T9� }��tvN��r�����V�����7�M)"�	�{�T��iI��}W˙�e�-^~Z�u���}�؄i�7dX���ܽ����d{�
��2�R�H��
�ʽ�_'xe�i���[�EwrbQ�^`���18�_i� A���9H6��?��}��$�`��q�@���C��#�:�E�|�+CאT�v,��#Ò�B5HĤ��Z�'���9��UK�<$<s�ds�g1��O�9Ar��s}]���n�2��X���k��O�Q�d�S9aNuQ�킊3��8���]g�U��8�ge=kM�LH�6���m�3�����9���Y�εH0s:��8B�h\|=�����(jX�=��� E�!j������Qe�O��c�׭ Y��	�8�\i$��.���\ �?"�l������F��6b��[7ۼt[y+�ڜ�+�