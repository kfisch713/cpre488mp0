XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� �;�C�s�o�a7�L��B�U���i�!��P��;v�p�B�]V��g�6�I����P������KN*�fP�
lܼFb�ʚ\tbw� ��G2j�L���dV7�4̂�ҥc�T�T��H��ޥ��m�ǝ�ǉa�2 Lg�[�%�H�?���r�����zcΉ뭺G�׬0R��*��Jܠ?{���#P�U(�f(�~�n*Dg��� 'M/Nt9�-,h��j�L*];����x9�&��J��H���D�䬡����#�C:V)B}��X�-�����"mwO� �6��>6�������/���i��b���X�`�c|�t&���)o�$z�҃�������O���&�'!�"�8����^+5c���aٱ�D2�X�,\#�܀91Э�2���kO���:U�	�Y��޳d_=I��,c��_驄 |N񔱜VB��sl���`M�{j tq:�fNV@�B���vs��88���ؠ�̶�sQ5Z���hW㯗8��U��Q�����ޱ	l�w��ێ��8��M=hse���\�]��Wu���Maپ.�{�h�~���	���S;_#Ф%�.{t����"|�f@%st����wcK0��T[�|W�X���x�YS��~�1 ��!�����i$c	(�*n欺e�;@+��>*�����̗N%H��q>rià��`�B�M� �s�dF��1�����"��]R�� H�;������io^�k;fk"#��ʳ� ��tXlxVHYEB    fa00    2040T�O�rFp#֧v/�#G�o��<:MT�n��=�����:�J��;ֱ�����2f^U֝�m�\,���u���m�����m8�����'�-����R�)2m�{l�Q�����v�������"���\�3��bH�SL`�A���uh��\�V��,�����Z@㡔�u2�M��ս�ާ�Ic�h9���u|A��ݭ�(�����䰲J`*��8�����#'�����U��x6���6RmX`ZM�� C-�i>"ayy�����x��!.R�ĳ_��
B�9�9 1�y��Gԝ��e�a�|%aq��7B�B����Y����C��!�Si��Q�N�����W���+�ժ��0����Kp���Dw�'�����=�CL��2Eˢ~�+6��҃���赌5�J@�];����@س2�W��nR{�v�6�$���q1͜��}M�<`
SXUx"�<��{CPSg��b��a�7̏t/�D!�C��i+�"]�NLg�֋�v������Y��:��tռ�� �-@Y����V�?J�`"wѪ��߀:A�Vٗ0tE�;���DL���k���al�&�te�~��S�Ũ[�B��(W��`����)�_��/�� �H�4s���(i20OA�Wv�IF����<�&�����g�9��"k��q�i/��:�P��D��׌�	� ��qJNCHvq�sL��x��셻�B| ��\���(�6 ��(���#���)YˌhBc^�4��1)�q=���� 0_�*�s���2�賭g��-`�E��o��O���g��"
y	v<aHDK%����wo�����^��g@�C�]���(F�VKI9.	��I[m^�J���=C�7g�ɹ~��,���5��i�	_w�L��[�XT��t�Yn�
�(��ì"�ψ	O4��g"p��E}:d�7���1Y�Ո�Q���2jfG���ċ �	(���}{ι,�Ǩrϓ�X��Q�źd�F��mb�=?���B��^���6žq�7A ugZ��r:��l�|)D���e��Z ����ۼU��@�:�t�8�R���}����W�z����a�w��پ�N*�6i�{=���������*�{�o�����yJLA�j�����*�#yOr{��#�n���Y:vD�i�\&z"���6�|[�s+�b\�����>�'�6�	�o�m�]ƣ�5#Hig���PK�g�y�%��`��q�_z�:҅F��k�ӡg}u��A�t����|����G'����B�g��_俴����2e���:z�wJ���Rk��W8���*ތN7e0���|#�ؗ-�ȇ��������0Eo�������>�[���3����ND� J���t��k�����ʹ'n�,&9 �-*͏8�o]��	ŪN�"����\�D��������Պ�c~�J3�|�,iҘ�c/�&�[ht|R{~Hw\q�3J����(�It�$b��g>xYӰ�Z���#Fх{%5
�x!�u�A-qL�����h�ä��e8eѻ���rt��2<.=]��r߲���	~���M�/~�� �Kd�Ӎ���U��?��nI�O썸��(�_�ϥ�����Zp��,h_ĺ�*�^u�YWXԂU��'a�qu��	�*;3< �>��0����5� p��US���C}�g�!�Q�����.<oG���A ?��[&G�{�#o�� �^a�煥�*���
�X�R���@�zl`��&�G�.-e�#�*!p�x�����ʅѠ�%�m�3�M%r����֕�zJ͐_�f%?��"�e4g�Q���Ý�tO�|.Ϯ��$�R�ď��t���Y�yl84*�;*r>+o�l�;:gx�sՔ��C�揟����qN'����xO��S�tf(����`DT�^�Q��!��*#ޅ�ÉkN�l�Z|y�+.�Hw���|l�	��7V:$B��p�T֋��O���ׯX�8
��`��=�o)�>F��zI2�O.�g�g�>�J)�v�9X�]�%" �$�Oc{�T�ˮ��!<fh�d25��
a��R�B���� xPa�;���E�vjE��.�Ƌ�#�(4�"M碪��l-_㦜����!Leh�}��;4[<�;��do����������!7��]��̊�@�s8�j�'���x��3u��k/2-K�+�i�գz8f�!C�q�CTQ¡�;&X�,��fx�L�c�TW��L���}g�w��w/���5$ ��P�j �5v�p��������ˠ��5j�U�5�Z؄ox(���%0��w���]�躴vl��bEܴ��鍣�"�F�4b�Nx��{;]}��ߺ� �־���-o%υ�vX���b���#R�*�;q ~\�elrQ 1�0oh����> �32��D�b�8�S�( �}=@���?�����
�Ֆ���H��p~�1C�2��CI)Y��oVx�V�jh�Q�-���3�����Y��������l)�V�ĪA	M��+�\�A��}D�h�L(�u�e ����{���a�kڄ�V7M�~��LR�P9MH;BV������ө��q�ٽ_��l�#2jrsv6���=U�!,�V=.�#z��@vt�'�VC��ȁ��~��=#�96�V�Y� � �ܫ�2�
m�$G'��Z�ё	���'��`�F���(���
7ehs�p��Nl%���7/�������\xA�"8�k��V��+7����w~g�^�wl��PDb�Z�9���FU׎���w���LI@��ksCJj��:��G>y��W�O��"��OtMп��e����[JvS=h�9�be�ݿuSk�¹��H���_���$�n�Ͳ+�x+b�@���4{��.���|Nj����!?C��śoO+Ӌ�&��f�d����Ï�Y�R����#Ӻu!�duǮ���eO<�Ǐ_��H�����u��7�i#���~)9��TGa�������3���»�g+��@EYz�4yߩ /wAv���M��_ ,��2�R�q2~Y<����<N��qs}(	bJP���@~�|x�P��o��<q.ڣ����/'p��?IМ[p��d�ȣ=^��,,@��-O������C�R}CU�� ���b+t����TE�7j�b4�6�-���m�[�\��`³��v���$��B��+�w�������qь8"��x(�Z�6��xy���䵥�B7�B�Lb�Qy���?�x��4���π
(�7����5`��yO2���
���ff*]E�+�����A�s?r(z���rܭ�4v�,�=�Ϯ]�$6�E����3��@-(ĉK�%���*uT���vZ���K�`1/Fl�?�K#��86�hHH/�s��{��v�u'9�L>�2C��Z�*(	��e�YKܛ�s3�00����4F;$��1]�S�6�Rz��C'P̛��>1�&h6��m+�z���}�a}�������
=8=�Ǖ��"��~E'@���G���hFvSB�I�L�ڄ�:�9Ԥ��@����6�Ob�u�ҷ�����,�����,��Їz����� �V�[ԍs�-[���2���2ݿ4����Vf}z�z4�Q����F��<}Gl�~~����4�,@+]�XQ?����;�G)�����mT!W���W�W�_9�g����*�ƙ4�NJ�RW1BHu�ŕ�xĬ��j�2����)�U��������i���1zZLw�7���^�I�� �@%�
�|Ӌ���v�'�f� ��Q Q�����7�i�f��]�kܰ��f�f{�9���p�6,����~>��_
$��5J��s�-N6v��7�7�>��	i��̓'Y%ݣ�a`�ȇ��2�%k�������'���Z�ۤ��|4!j�(��B�YQ:�v��/7[������y������`;�tw|��[��Duw4�����i	K~�N��*c����E��N�p[_�@��Dõ�����[��^��;`��H�G���6)\ ٯ��V��Wo ��gN�H`��6�k����.����Bu;��ٿ��S�b~������Ȅ��ӑ�*xεq�d��p��Y[���Nz��ۣ��zb�z�Vcqfϫ�4J��=������Xg�L7K��^cf���g�帹�}�l�+�È$At	�$8�ֹ�����Z&�u���Q���G�\��Ӭ�P�!��$���ł�(4#�[�P�퉾��%u��t����N��} }��a$XJ���oB޽e��X6L��α����0�Fn��Ո��Ogx�jx ��'e;�n�(��YT@�:����+3z+z~��<8�}�%��׀�q��I�+!�$�`Yܯ/�U�y=���j� g��X��*Vkm�7�w�0V���\W
�G ��Z��=�����O��{��Wxy1�4���;Sb���r�1��
�!�~�R�������Su���Tݘԑ%��]�$-؜kv��/���Y�|�W�M���A��=�z�)�L��0��:ms,�:
 5Pe������=CfL`g���z��{0,����o����g?wv�E��U�zЏ���t�$:�K	e�~Em�S�
�ފq�!��q�4I�����jM�:Dy��Hx6o2�����QE��Ƈ�q���?���	�HQ�u�:a���
��*I#W 9�����-����=��Td����E�8T�týd?�W���s�]��{��Y�V��� �ҷSw5�u ��(�3}�����i�����=�0�1�$���RH�:�0S��`y��)�}[���
�н'Lr!�\��G./�SaP����E?V�ߴ�v&R�� \���"o�vT���z���wڤ��&L�@Q��g�V�Ėv,��f̶F�vI��%\�F�,�:��^ݎ�1������S�87qt����ps�����?Z%'=��'��+��D�3��e�����O\�-�R���k�gb��)N��-�չUdU�j���q�����t�j-�]�j�G���C!�댇G��t�
�_M�ι�NQOp���THP��h�^��l-����Ӏt�����Er|�CԠp���L��[�a�'gNR��IM���qX1i���ʾ�b�Qw�ܛ�w췒�����t��f�1I��V�x�(�\�XP#1�璍�[Ϛs���Vm�`�}Z�:�<�ȧ�\�A'D�D�3�7�:�X��n �W��'_/�^n3���:�:����V^��&��z�{��Oc��7��se�Ε�K�~��p�r���|U/�P��
����lj��G�����C�}�@\��t0qV���X�{߼0,�q�,G	ށŷ�sY�Gp�w�`�������[����Zgvy qV�E@�+��Tf�2*��K>�*L�^2i<�Q� [&vf��uޫa�D`?��o�x�E�9�O���[b��qu,�3*^����nT*w�FaV#E�$F�Gt�Җ�� ��oL�a�3�8�o�m'��r-�U*LSG��@	�!K4�w���:k��Z����v˝/CE*Vֳ'�:��mAZ;��_�[���(���n+G�F�+�bG��,�;U/���V�M�膉՟4<�������Zv�s�(�Ӣ$kƮ���@�]�6ƙ�~�2��n���j24S9"���9�I���Wաly��Ѳ3�®/X �=�(�^8b�g+��Jn��܉����eR�$Ҷ�O��
��SAsx����"+NMA�id�[!]G����R@��e��+��<G���C'{Vm���r���"}M�;���;��y�|s�C�~ !��A��/�^���FҰ;l�	�����������r`:"733b~=Ɗ�t���P(w���B��A��kL<�\�y�v������� 52�2��|ud,5��oN/zv%�M�W|w�қ�y��ؒ����Y�\1�O%=��5����0�<�k��ѩ�ƨs9�z<��(�2���hp�����$�<����i�	�.�S*|qP�m^be^h���e��@1g�U��2�Y* ��K�ܘE�ͪ�����e-�����Dz���]���[	���;g1 ,������h^Ӵ,�[<�]�����V(���2��v#r�A�ߢ|@�~�����~���B��͓���H�Vx�.��)|���W�¸C�n�$PB�}]�Yog<������Ĵ�/B{��bZt9u��d�/*�ӋY��{+B��_�d�Obb��n?�S'yLi��G^���H;;���?J���3�>��t�8o�;U�' ��	sU�9پ���t��WLY�?�5��b����;S�'
{��O�����	��=�)\��!��ܴ�1�k�گ���"��I�n2M_lf(,x�}(���'�]����0E�����K�Р��DtW^��΋�35�E�ܝ�#}�}B��z�H��(S���F/ox_/�6~�L�k�+<V��0{j��B���G_�Fk�-�B�y&-������H���u1Ms
����	���N�m��&N�V��[�7�9�`~����F�[:�@��K�[K8����S�#�^v��?���+R��d�ú�!������p��8
��h](Y�����AF|�O	�s>����~����ȼv�b�o���4"***�"���� �h�T��dP�6�:#[�͎����+U��%�;�Jo�%���\�.b���j0@�H0�J�%���à�~�S.��[lJP_sB��iݠ!ٿ�3�~�"�Bp(e����J,�H���b=e_��N�8�ir/���?�wJ��:�*��LSZ?���8�����������@lE�l���98�LCd͍��_�v�.>#��+ �r��^S�4��L>�߷{3��/��e_DM�z��d���rS�]�lI���ݨ����=����ã���u>�=3Sn��a��˅*Y��ף�a%�N���ɂ	b��ݦi�n�e���[�1�Z�t�y��k4f��S��2����L�m^qrӺȾ�ހ��~L��=�� �D��GY�|���m��H�i��V�	r�k�a���O1���fs���~���֢�zP����jo� a�(�@Y�t��C`��TP�m�Ĕ&h8^hZ%����\�t+a������p�a����(7L�}7v��5g��	��,�v�=.ÃW��=�hK����B�~�iI�ج���i��o�
��G_��W�Q���]�L��Uf�����5%���`[xCM���NrV���������VT�L�8pxy����-�^�*z�F�faq��r|=\E��MV ��8��藢�����rɨ=�GX�<�Ԫڑ|F7������������sвR'-�ʴ>	=�F��~Y|`?������}%j��.�'�������Jvg�D%Χ��2b|+��Q8ޣ���E�����pZ�E�=kU@�U�ZE����<�8���ة��__F Bxw��q����#��
�in�Ӈ@��l����&�MO��N���G�m�5�/��M���H;�;;5���7�?q��|P
8��������D;|st�p����n�����U�-��|���Ix* ���n�C�j%�<<A/7��
�͞bF�e��Z+]�_���zI�4�~�7.&$�
 ����c�S-S[u^:`�X��өr�����[͑
D�~$Ԩe�3p>���6t
Er��7X>�Z�|+��*H,Y��{�7}�
J��kMA���f������'�Y�z�y����n}��u "v��is��K#%�u���9���M��\}mRb�m^;J8��<��g�~M)���d�ښ�k��r���#vЃT��I����a��-��'��8{�Be�Z���ꗮ�
m����AY���Gmx=ga�e �l\��a��m3�W���#�|�A (n�$)�~�� ��W<���s"�8�?�YQZ�	�8r�>��t`�WIv�k:�G7H�c�/������6�$ù2����ISFs�%�X:0B�D
�PX��5�b�zS�E���	t�[}L���a�呄:u�B��FM�̚��%\��Z}1���,���RN�l��E��CM�ؽV��L��tN���S�Y3w��G��c��0XlxVHYEB    4f62     b50��|���g���Z�Il�Yl��b�����;���S��ސ�c�2b+���ś�'=�hȠ���٨��/�F�_m�Qe_��ŕ���hN�[zQ���!0��F4���"t�o�����A�>�������%1�`����=9tIxU�kL�i���S�uB��V��jɖ���皥�<�K����?&%�w��I5F���)���`gr5��ҙKc��8竈�3�O�M�4���4Jd� ��[1r�x1_� ��1���-�`S��O}C�w�ʰ����GR��[=ޝH  ;��J��p|�ӡ�̡.�`蘑������� ">>J9�p.F�T�q��u�����9+�2���mE��N���\U�K��1{ch�t)�����a����3%k&׽��}o����_���:�"��N���׎�]K.w�gth�ck�h�v؝�����lh��H������vn��J�dY���E"8�vu��##��dY�E��Ƣ�r�,j��_ݴ�=7X�J6=Z��ԭ�N�u?�S�s���rQ�� ˺V��k�ʪg)�d�bE����!ƥ�|pnP���ʔ� ������j��WU�=ٖ��3U<I�~���^����?}�� �'L0�5�e:�-wÉv�f�`J��$JD�݇��\�Oݕ�z�ί�-�]ѝ01,����-��O��.��	$~P��l�Al�³�*���^hw��ų)p�T��&�a��}�W��?�ߋev���|�@���8*����pL?���3/� ��QB���ܬ8�W��,��̧���O-	}0K2�Κ��%�X����{�<�?pY�J?�18m��ɫA��Åg�1.
��h{]o�r-�!�;��g��Dl&J|c�Y*X��,����3`� ��t�d���a�G�����x��
9-ΈY�|�9�r`V�wމc�����
nAB�D}��S;�"��Ƕ� H�����ƫ!T���
�0'���<��w���.t(Ew��H��5�F�
T>X�~�V�� n�!=��l[�U����0կD�i)2�<�W������)�n9Z� �4�"~eQè��*�?ꒌ�6�E�߽����Z$btt�x:8dB� �ű)��q&I���+]��-k&� ��4���6f�tD�Q���Dz��zW%�O�P��'��,=2K���l�O{혧��S4S˓zk��'_��|��T���4��4�����]��̟E�P�<JP�EM��\�@���k�Ɲj��p���T3�_eUl	�B1�N�2�nM�2;\����T���<�`����>�0�x����c��93�v�H`u}ړ��V� �>�r�q��rW�%�f�
*R-�&������
T�ѧ	*I<�k��t��ܽyʂs��S�|'+���߲d���c�F��pVs����)���T�|�6�&h~�p��=˞����$^��S��*-�a%�s�vuu���p��}7\��4�	Մ�&�iܯq��q��IVʨMK10�V��9�m��rcFr5�Y���c�5z�hm�pv �'����7�A�\D,�vR�U�`�iH�zc����LJ|�+6�⿵�]^��r�`�=^��	XV���2J�b���Y�"2��87�b���'6/�Y�ҫ�p��K�y���k�) ��9�h���X��d�i�\
��<W�ڬ(����1l�[���f�mw&�M�JM����%�O�O��v�+<�?�b��B7`[C#�k|x������D'i��y��ޛ+U���	��ƇT�ΕqD�S�썓e��AM�Az�^�����1΂�mU�qBa���m4��?��'��F�+Q���)�?�6�{�e�
�A?���IXV���	:A��������5��e�p��Y��I��e!tpV{ r��g+�1��6}�h�Dہ��U���js	���`-��N�}��)=�����3������Ƴ�Ӗ
u�
�cn%��a깻��aW����4bx�7���(�W�oR��I.�)��:���wsOtZ���'ɰ�Q7S~���g9�p�RD�����/L��+�U�1p� 3F����Z?�ʵ�,��`q�'68O�eP�:���h(�g�1��nVК��b2@����|��z÷v�=�Hn��xmTi�0Ϩ�g:�MN��fB��B60�SGz_)����b����!`�ַ:D��XLH���m��M��҇<k��\-����l�ݿ��"+mfv�L�rRj90bvh��܀�)j[�A�5�R��ʼ���ԜHߧ������,�%�|6z�:�~�%�6{�|�����A�w�G�w��y)L�<�μg����%[2���+B�؀�^	���0r�E���c��"f���iw� �.���/%"t�������݂78@��&�!�����l��h�G��� t�e��!&AS��Sr.�%,q��E�..X���R	`�mwy���} <xk��%)����I4F\GRح/p�xnF��o�f�%ϸ�4��"H���-�Y���.Y5�+����R�k����}~)r1�K�d�-�I����Ș��U��Α\�w���.ҡ������+?�rYa ��Ơ�k��O�¥Z[�i6���O�5�n�DZa|�#��q`�H�飤�ѥ��aa�3X׈ b�?u�THX§�]��6t��&��Hg~��MuJI�c�qz~O�<xF�5p��,�R�]��9$�q�B�@��a&�o�P��cN�#n���R4~?)�F�Oǁ�e�YK(�{�-ʇw����J�3�C9��	����P\P�f!�,���XL�J���N��~b�(P�e\Hۂ(~M-��E��n�rJ�v��(Ү	A��P�x�S �J