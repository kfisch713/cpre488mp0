XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0�Q�߳a_F���XXE��%bcBrׇ�p�a~�E���&��|%'3��_�ho�&��;��TM����
��(�>�����g�'䊺8�T�>�s�����	�q�h�S=8G�S4��
�h��y�l�[:�&���vaf:+)G_'�#����"X��N�ع`'3�\}-��i�;_p�����fC��y�>'��y�4�Z0qU���0:��<6>]��E��/�֌ݝ���9V$���%����@<�!�(T��'Dr_�� �-�f2w�⢺�7*����5#:�&k���Ũ��8�6(#t������l�3��EA�)} n�Z�;k5��q#vx[����[w럹��8r|_�2����	)���ҩj6�p���YOE�?@�Mz�L�ë\�� ���UΗ��{��nYs���)$'9��x�o��^�
��2�"<�j��8Jq��V����w=D`��ެ>Ŭ��#�d����*��k��8��IR�\=�ɽ��K�-�Hu�o���NK�b�8h���	����[�:�������0*>�PU����({�WdZKs؉m��;:]�v(���~���=�a���6�
��jHɠ��J��8Җ%����p���;c�WsTOl]`��܎��E -nb�U�C�~"�)�M,0q���bii���O���܌<�gP*���YG)J����B	�S��Y�?�ʧ��H��!h|z�vh�7o�l�޷�}c�*Z���&�XlxVHYEB    6014    1840K�_k7��{�a~r�~�-�gRkc�bwZyYl^ϳ+�J<�x�/=��ktІ�?-�n�8T�IP� %fn~�R���k��HjAd��r��R"��G
|$��W��(q��.
�h�T֑nU'n�=FP3�h���􊖀�A�G��� /����ob6u����<�+@w��j|B�Ђ
�P}�k����m���n?ə�嗅q�x��*;���N����[�/B��c
$�!;o�Xx�P@A���������V!��|)؞��җ:�`��O��d���t ��1��T#Ek�4���V'M�� �	�8�ʅ���jR-#s]�����Kh�Q���A�1�i��iO]I�`��ɖ���Z����N�D��#�4�x�+9��>D9��t�5{	����|fV���[8�\���A�x�}��<������aI\!�z����J�tQ���ȑ<L���
��΍��x�htND����-%��-A6孡�D"�8���s�'�=�	q���pi �c~�������-�������'V+�*|����>�UQ���_Y�6sp�Q'��������$�`��.�ɲS�_��a��zƽQO{=�]����hH�R��}|�)����J�V�r��Z�-�J��Q�c|��1���ɓ�,���q���q�)|��n��X_�OGt�	C?T�d��%4l�k�!-ɊjO�ʋz\6{xH`�ؗW�����Ի���~;a�71F�h�Zfe�%�b�u��,H����SC<���*K�Q��+[���hd��I4K�E�Z~�z�{��{vN�HFp���r���+b4��}N�S��yL�zA�c�����w���P2�Ӝ��wq�
CH���e�zǌ���5���q�h�4Ю\} �&#�У�×��\S^����Jk�g�5� ���ߒ�t�{�b���^���}�珠嶤@&� ����bc;%��+EW���B���\������;JW͈��¢5���(����'~4�5We.�}�ؾ��=�3�Uo*��g��D���UNm6+�Z�яM�Pg��A4ƞ�:1˟�&t3�W��b�����5�E���=����TB	Jl����mM�m}�;{�Q�
Y�5l����;?��yc.}F@fq��xK
�Y$h�4$Ye,ЄMj+(�C����_V������K�s�>��<�����~�L�t��r�0貥�}AH�Tۣ �-P`�&�j�ibOa �
�;&DŢxc	�Q��\� �����D9O�����np{[���Rl�� ���XW~e���*�O1�wQN�6�#jt�+-� N��a��(tQ���#�En��_��C�/���A�qUT�9��;�{�Ƙ�\��&xL�K�z	�IbO�RI����-}h?���w��hnI��C(�;���F�G�7Uì!��f��9�P�h���o>�z���?q&�H�R���/-������u�hmi ����k����#���_�U��p.¾�ީ���)x���vpܴ,���A�^a�-a�	l�F�)Y�yb��D�v݁jR�d�!+�N�\�n�ɒC�������L�ƽh���\:�i��U� Ԗ�=<�y����6��<�T+c�큻�C%�nj�&o�CU	,���V/|J�Ac�\,�l����G�lY� z�LM�U#Zv.�P$���;�,W�������t]}�@�@�j߱]<��C�Ԯ�Z��o?�ĭ-�����p�Z�i�;؆:3�7�1\��1�9�p�{�
��M� Ljbց5^!o���$��{
��x�`軙3J܄�''��x�e,��X�E��^�q"t'��qf43����d��.O��z#To� �&���n˱98�w�
t:y�-���[�X��[�1|�x}PINC�Z~�f�A���1%���
�D�*R���r�sܼ�H�@����0[jL��pLè�������p��z�qp,~[�3�ķ*�
�TQ�6jh����^d�޾�k�!�v?YI��ސ�1��CDTmc�r᫩/���F��lJK�#�f�a�
�J��.�)f�*�SQ��p·VMh���a�Z$�[BՅ��t�qsZ���u���	[��q��¡6��'��=�L��Q�����X��*�@Dx�ډ�ť�ܰ~�Y}��N�	��ԭ3L����NO�P9n )TWa�^X �,pH-�ֲ���t�s�3�8���ϭ�^����zY-�	Rp\������j_���_���|��r�jfñ�	����\z�H�i�}U�0��Y��3�d���u�8}�f�iPG����}"��c�Zy�yj��;P�q͏�	kT�5�k���?���y�˫}�ڍyn4�d�Y�G/0����_��%���ɯ���z��Įܕ( �=�f_��|a�:�m(*��iЉ���57rj}3���#;1�;�6?��-2$M��΍7K�X�({�J��<m��I�[��+��3���=��	/��9�P����1�Z3EE�TaO�zG�t���v��ԝ�L�ߢ"/j@�7���5����>)�r�!�� i�i�T2ɪf Ȗ���#��2�|'ێ.�~tfr�~s�J\��Pר!&	� �G�1�y��pxx���"��a��-DZb�a^��.2!�9Io�"5����^�vqONv�`�g%�ݧb���{�P���ٲ㡆އ�R�f�	9��]���]��=�����ְ�V{n����n{N�z2��9��O�p�{O���������Z5ٶ�)�6?g}�
���#��Ԃ�	wLp#6�1��,T��U���F�?�ƀ�ho��ݺ��e�:n����
%{�d�s��B��Y�Q�p��qn���H�	����%�7N��=}"����ش�?�u�W�GY|��t�{�8.����>��g�Y��{�����R#�$��H��a��Z���
<_�!��S�"�i��T㩒���d`<��s�%��Xx8{0�����@�s@V�x ��XsYuМ���H�1��e�\]�\�a�u� ����9O=����؛D�W����*@B��qϻCɬ|"�x��M�2p��LQV����/��|}��e����������b�XgqƼ�f;Dj�Re��5b����c��",�H_�����y=�Āy��J�%:�C�O�on�L����R, �^�S���<�=�#2S�01�M�h�Ⱦ]n0G�����t����^�̖��:?|�_s݉���I[9����L��b���c�Y�e���2��z2m�1��9��֥�0��&�b\�Br���d�RM�%īrUx�Q��&_>|�N)��}+��5d3�N
.B��JFU�pc��&o={͒�2�����3]	Xh�����S����kc�|_�ǘ�I٢l̿$��ɂG�\��7��v����@�*9j���݀j M�[q�JN�G9�g�]NZzph9�gAzv���\e���SV�l�B[�׍�D#g���Vj@��z}�r��Ƞ�X3�F�y9I��4�/����UCg7��M�,Y��+��ש���c�y1 �����|��ަ�0�_��.1|�^o})��9
�Ebŝ�b�a��6[&W��
�z�ƾ�aB����u4A&�h�˱����?�QS�V�R���!w���v�Mm��u�~���e�Y�Ƚ��Ӡ�1 �Q�;#��~�Y�\xK����s/���7��r>i~_��9o,tx�-\	6jo
��I��+jF�������cȘA0EG7�ט��,q����-5���L�0*�+�j����9�4<���Ҡ���=l�q�^N���3٠�N�bӹX,唃[켉�$ԽXc-/0F�y.�d7Ȑ��1Ls���D�j����ӆ�<�oe$t�6Ϳ����6����5>!8�����!���A5�w��)b�_�o��m��n�͟�)�-pG+}eѾ$�[w���1�~,3b����Q��+���Ee�A7.�m$�D��	�~�.7� a��������,ٔC]H��y(�36���-�	ШnO��%[��EA�Rܛ��OG�o�%+��6]�T%�NyE|/(`)����݆�?g#�LO9�S_98Io�gK�DG�,��ȿ�d�l�W��
J]�z%F��\9��F9��_�h߱�W����-�8�\k�п>0����d�B+��ʝ����R�����Z(1�m�Ȅ	��R��^��D="���S�]B@ض@��ӹ�{��M��a5��B[���LK眧�����\B��㌿�!7����u^:�p��'=�|��:�ܫ%eS��[�Q~��'��P֋=p��~�yк�w� �T��d��������^fIv%���h]�*�"ب�Y�C�*�׍[`�5�� �6-�Ri|��U���&��׭�ټdC�b�G}�;"���;!h�-�{
0��2�]�_�6��/��ڼ�cI^}��ȘP��c6�'G'�(�ev����N�րB�������e�Ӝ��H�u>���[���ע�Y}-Y���'f�����BI�f��ȳB��vMT����oYh8��Z�?fR�G7�k/��q��y(aP�֍���KwwA㗈��a&�!o�	��ُ�C޻̦ղ+%�4��s�7-�E��畉����)+��m��Z*�e ��xS�Zިc7�c=.d7�{AF�i��=�a� jz�*O��vO6E*]+�[DB�*�QhP�1��-QRHFQ-��+�H���	 �ԩ`0���I֥O�´o�ZAh��$ ������5�O�;n��en���-^�ΣJ�Eښ��G��F(ɏh{���@y�������EvM.�������4qu�z��d�ql���f��rЭ\X�C��NuTkjP�2�i����ZefZϨ*�v�#�U)Hc�V�Z�J�4�ߕ��o/?f�8�TT)*ON>��R���ņ�U;A��{�-�#�O��h��v�f�0驮���~���KM�CB�O���e���C�La_t<�\'��-�`D�Wmv���f[���yy��bh,/�|�A0�cH�(Zs�*Z3�r��?�l���(L���Ȗ2�XRRø�z%\��G�1;�C����N�����|O�o�.������A!�}f������A�k�C!�:h�>���^ȁe��M��8h�c]�����♐��U�N%B΢�ȓN�ajXx�C�9n���(�D�E���@��t�<�;���Q���v[���=[.R�Z:�<+�5~/��s�b^a^����H���#���jHc���S*F=�sLx �N��]�l�م�7���v����a^J`��,琧�Ilœ�#�snQ$�lU��\O����Q���?�GP[H����i�YXYi��p��["%��w�����E�x4vSܪ.��$ '�:����3����
�(�� '{�P.;IV�ɤh��g̜n��.�-��$X�1OL�� 7 Yz��VB��ޖ�s��N��X�����e��SB�<��x�lSc�*	~���L�_o�/⽼r��!�
1Q��'�-8�y�d�&�hK2STcs��-�`ʡj� � 4���%�9���Ֆ����q�B��n����e�?w�ffJ���ꋱ0n��D�̀��qi!_�,��s��ա	>�6��I?5�2;�Dޫ�M���c��W5���"ٷM�W � ^8I�I�8� �о�z�9,S�������*ɕ�Rp1B�r�="�Ж��$���r]���HA�
̴�(���)eXDd�-�=���Nt°Pv-�G�Hq(�}Ԑ~��4m��Q����_<� VH�A� ���r�61�8��1��B�X�?�k��~��|S<�&�3y}�^J;�X1��Rb0X~���׀�~��fP��-��~��(m�8N%|�8Df�ʷ2�$���Oi��K���C�|o`qN�^�K_�|܎:��{��q1�4�_6�d�i�/��AY��8�C�b���&����c�8.?c�W��dn�.*�A.V4��{o[�������x�������4GƑ�������{�0��ӜX��Sh��C��K$_��-&��z���K�A��C�@P�r?'!2���P������y����(�%�