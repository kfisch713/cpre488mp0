XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��]��Ps�o���$�\���5�r�+� �l.<��%G<�7��d�R0+� �4��R����?5��c�lv�:�3��!��0c6>�� ����s;�0�X'��-u����Jg�%�� ����^d�T��J0T����h��jz#3%��Z�&A�c��}��!��)�V�b��Ͷu#�j^�1��jt?�c�ȣp��sw��s�&9�����7@�h?�)5b��_
���˝��#=�[\R6��}��K*�)#VxX>���ܟ������d�#?�ЙT�f�"���>y(�$I�kNʹɾyY40���}��/�Ɏ�X�(lG
�n�y���q�+�%��M����Gk�amj�cmp��ǞȡԨ�@4���K��M��7��1�ի?B�m#h)xh���3�0�h����a�Y��%���z��1*���1
k����ߙ&Q�C�+�{�|h͡󜜣��'cd�1�`qn��r�)"bm!h�v��'K�xG�x7����t�J�,$��t>N)������$�״���q�U�[����/˩f�Dܭ�	I�[�i��aZ�5Y�.xio����g���F_MW���yah<�a@��dK��TV9<;��E45������8`;��K�gM� �����T�>�"�0���|$�����t�`ڼ^pQ�����?�l�+�a�h��xoQ�p�H�RzX�j���j)$�}a6sd�1�j��y��WW��n7`��㣖���r5m��2��s�@@�D>�VO�	�V:h�%XlxVHYEB    dd8f    2160�_�B��g�s
C֞=���'��S����]�fJeFS��K��#`7����gl�-͗��&�/]�Y>?���%�<��&W��5U8ˣ�*]�)=�-i�ܗf�Ϻ?4��Q&.9r��+�>
a��a���(�`��rO��u),v�Hݦ��V/7���6f^��p|����~2�6tb�/�+]����Q�r沝���_Ppw��|~����dX��"���n7�D����#E	���憃��"���ؿ�b
`mO�
n�Vae�L��t�b�VmՌ�^\���L��V[HYt��=� 6r��b���ɒ����d��+0_�Ս��F p@F,&�(۵�w���6F�7�6��=#�m�uyk�n��6��[$��� �4�@�~��[Q�8M�=X�ί��H���%�g��>���XU��R	�/� 5$���x�c��{��dv&��W@D��'WXk�������#�s��6S�R�;��$����@��`Y����8%]Z� 3H��j�����9'UoLpǺ�y':F��^�p� �R~��4p}� ��������T�O#$Eһ��+�i���Hv�6L�"�#^���ۢ�ݡ4/�&���-՟�W����L���a���ė�ݐ�Ө��dv�H�~%��S�w��h��7r��ؾ~eA�����ً[W��t"$�]�sl��f,���������w��Ҙ3��;h(tN��jO�*/�я;�&_x*��/J
�Ԇy*�L#�6�s˾�.�20կ�2�蔵֧}�� t�QѢ��"Il�kb[.����I�#��<�y���Ł�\�(�&r���.�1]�(�:(�-�r.����u�<��1���-�	�os���ԏ�.��oR���qO��x9�*�Aiʡv�;�{w;��`eYG�?��*�����#yT��(�#x���7�֯�BЉI!ɬ����ϊ,��Fr,�Zѥ�����m� ����fuf#&�ɻM�p�VP����Έܷ??��m*�N�����U�o]<����YSz>�����V����$�Ͻ�Wa��z���)�|�*�b�;���=�J�5���{:�{[:�c��x�:@�!�Mg��s�������a퀮��H�m�:龗\��;�?�%�V���̋��B�ە=s����~�)o�?x��%N�� ;)j�yHŌ�E�.$>�|{�(�.�c��,���*� .���SP��%4CVSTiJ)z����P)t:�`�ݖ��:�U�j����_�S���_��n^��.@5鬸��ɿ$�W��b5�)�`s�]!��I���u�rԆ�އ��"���7�fAo��^�MŁ�ya������M��rR#7*�����`xC��j���ø�q��hy�,/�ߏ��G�4��* V�� 'ˈ���N��+����W����Hg�G��6��f��:��\�?M�P�
͝	H+�7-x��Q�Qq�D����"���n�@� �6��y�l5h��ONP�\WJTߒ��R�H�̎!�=_��~����-"�4\ �i8p���L+��5�Q��l��S������:�SH�ɝk�	���Z�m�U�SSB5�(=$��]aV��lsN�~��T,~��M��&���@�=g8F���ic�ك��+����/� ����nƹ�1?�����n���&)����% ^,�UV�A�r�����ӊ��.ʜ�u1�}6�%	�vD�mי��oe8@�S]�p�̓�hx�2�/(cئ�O-��~u���Hư��dB�*w���X��;����s�P���aw�C�;���c����E �H�<� <v�̜-:8���+�1[B8�A���c���#U�5��}��.��N�k`=�A�9���S�PoI�c��5|~�Z>E�,$�y��y9K"�Vt"6K{@J�9i'U��d�Utt�Z���(ms^]�\�,<��Y2){�?��Xw�|Z�a����D{��F�P}��_����}��J�}�-3
���k��#Y�Q*�Ю�e����5ʤF�ASJ�a|2��i��ql�O�E���J�3�k�y�p��{�Cs���-y�Ǚ�j���4Z��؉ցU�5��!w$b�>��XT���s�F�ʹK���W��.�G��b��d��ա"P"�H������J�߰g��Kkw�.�ؚ>��!fb	M�[��7@����|�<˰@�6��z`\O���q�f��1�H-P��O���|O�T�;�cvx!�C�_��o���g[�x��TA�L
��I�
�*��4V_�X(ڰ��[��^�~�1SD-������Ȝ���/����n���b��^��+���Vֈ��*�ë�P��
Qߘ��}J���vb�N�<z�����B�����ϸ�B�WH�܋AL��C�iK�E��<
�醳0�>����g�γa�!窴�st��K�Z~uJm�!�(�����y�sT�n�Z�0�����̆WX�`���'W�N=�&R^?I�5���m��K�Z��!	�\���e�`k�ؘ��9�>�V1�5|!�f� �n�\Xb�[MΚ$\QТ^!�D���ՄJ�����YJλ��h�M�z�~�d����%6������.WB&��p�s�@�X�A���3������6���c`�XG�EYq�RNC�H2т>� ����z���!4�
�spŊ���"�;Yh�� {X�\<|`����kD1%�A��Ԉ��7���)���M��vշ��$ěx8�&(�Naȍ2��f���Dd���GZ�� �dF_��\�p6�40,�9���Thk��S���[��zCQ�h����S"E�46- �E���R~���Ԏ�=�,j�x^u�I`j��hi�������������>VC-%���`X�!cO1�����ZJh O�\:6���Ds;6s.��,x��
����oǧL|���� ���(V�u�[M�B묧��0t�\b_֝H���!Ǚ��n��&�ZK�������P�,�4�xz�cP�_��ǅ]�r��H�,£����c��C����^�iro�Ǩgr����(�8�+\/��B��c~�h�g-��]�c��'7�-��`���#��Y>��N��ɨͳU�����rA�4�i�i�<L秥�H�Yz��E^`_7e��s�\�ss(�� ��O%�U��9�g�R��1�����EE����x
���X��P!���
�\%b�s�)1`d��?F��5&ݖH�9N;���-���g|��1�I��n"c�;�}�7�3�A;b�-_���P�:l�pGG��c[7��9�a�X��y�8�#�E���ڿ�u�B ��ܩ"�{pfLI
�����p�nz(��œڇ@��?����R;��D�.U��qac����a�3��-"=���U�-��Q����yGT���]Ŋ�P� ��N�W!f�M��Z� �ɾ� M;�Ŝ��B��RC�$w��a�Ϫ0{���`R�kj��!#�}U�Ty�o7c��m
�<Y%�z��˪%c>6��Y��0!T"Ϛ^O��{�y4k��wRk4/�u<�
u�P�T��^��N��1uH�}/i6:{]�r�����xWۣw1��l���ڏ��[e���ؘ�7c%Z�$X9<�g�`y�[�5�h�JH��-L������O�ʤv&�~�$0t�R?㡭�ʇ�r�f�#lI�1��V�5�j�����C[���ʞr���Ŵz���"k&v�|��ND�����1! ؃T�b���LKådw��g���=�Q�ƫ��O�+�����6��M����Z��5�� ��:m/�u}�>;q�>���5m�aX�'��ǚۨ�c���b�QxR�����`����,Z?K{���>�[賠��=�ݟ��2��w�4%>�E"gӪ�weBP��A�@��N��*Fߒ����e����~|ܜ���k�U�I����d5A�Q����-�5�R�P>�u�L]����n؍ǊC�p��:��+y=l��A��^JTB�Ir) 2�+���!���X��&�B�8_��y*�'����.�����s�c��M��4�!D""r�4�@3�s��-��� Y�n��PK��'F���[�I�
ʕ�6f�G�@F�����-uĄ���
�k��Ϛϓ�<)M�C��t����W;k�
�'�ˮO3��Wc�������5�_6
~"�!�m�k�k?��|��j���'���4�E@��n"U��h�kɢ��M���z�����P���j�s��B�Ts���S�V}T8��F��[����=�D47�wL�ǲ����'�_��G�D��0D(������a[�W\��ǞA�졌�ĮM�;�[r�-��>�2���!JBM\>|�skd�w�~"����^	��cF!������;���'�߆ʕ�ѱ�K�t&�R ~T�((#�.[t�[�Mw�og�� 1�pF�3�U���ϴ�Ű��8�*mC=��Z���c���L'sJ�Pɮ�CLx�(x���t���Jr �Z>�����T{�=J��-����c��x�]��ʴٮ���6� ��\J��p��N�G/ݥj���.@�2/iU�+b��ή�����cBfk�*�=��m��p{6�����v��~�JZ���{w��e��ˌtdeoQG'��f�d_�C�����q�d>
���k(%8l3M\�����U��z�� �Fc#����O$m��"@�]���߰LW��>����]|f&�lD+�d������V(t� ����tV|������'�U �����X��A��S���d����WcW0%<qS'��F���}e��0���H �~9����Q�O��eu�s��*c).jC�&�W=�Ȁ>�.�~8dgI㛴Ǫ߇��ڠ^�߻z�����=" ��< ׅ\��9����'�ʈ�GD�����iT��{r<�˰*�;�ZbӁ���@!��
R�� E�F�h��K�a�P�u"�ܧ������f�����^�>�$���ߺJ�Q��dGz
���e�	�=N�[ӳ�h��%PŏK&^��=�֝�k\Y#�DkQ*3�U3��op��M*d����Dt7q� �*�>���3v_��.��a =��u���C���-��U-�K�5T��pR��=�	�o����5�y&N�	[��،��B��7SkZ ��SID��NX6���I5�(�C�.��� ��=G(ƾ���`cM�̈<�O�l�@-��
2ͳ3뱒T��~Q&������O0�x�I�I�y���c�4�dͪ�����۱�����h 9���)A�w1���&n�p�IA|�g��!�Rt��*�@��Z�գ��A"b��\�$} �7�0�;tj�֔�o�36L }c��WÅ\�gz"���R�C�*E�Z��^��O��	q��{:��G�A[C<�Z�1�m<Z�,�K�Gp����p�'u~�jhd�T`�y��I��/(,��IYt�p�*��&~Z��2��Kfۼ�����i>���V������Y���;��(	9���欥��J煌��;) [G�@����u���}���=�]�g�������9��dF�i0Ws���s��[����;ej���K�hg~dѦb����5e����#7��#	#"CJ�3j�I:�6���K���>��sp'U����)��[rVv��{ID���k�Z�\�2�oǬ��yn ��
��wEH�_���&O�c��(�'�cj|!5/fk~I�f&6���fO�+�pCsK �8j���OpPB�V�i���p��C2E�Idt�:�O�
�_U͖"��������^O*�+�VT+h�V{�1�Ə>9&�u��>�,{�J�i�'x���:]j�"���H-���I�*Ec�!m�;y���lg�6`��#)҃�a�HtY���8�!jX�yݍ@G��8�Y%P�ÙTG4�$D���p �������+����'o����y%=S|z_����/���@��3��#��L!�9���hi@����K�g���/��L���h�^2����o{,��Bz}�1�#�P��n[_p���֑�c 	��S���X0���g�aZ�!�	Q����6����z�Z�}��+�+��J5.������4��sj�Oc�sRc���� �(�(�O��މ#���N/�$��*9�%�Zm�z��TçY���y�C��s���܏s]z�jn��gdྙO�oN�ɧ��wL�x{7 �X�tT��&|��0=��Wq@�45cc���]�x��>?j���/D��C.����C��2,1��r����B��Vۯ�%_���G'g������kk�J�u~/�:5b���i���]S1`b����{�+����e�>>&�Ym�r�oĂ�l�3���R\m�֤w|������hë'I�_ET3������h�%�+�"�[4�6�}y
}7{V_��O�`$��w27o��F��ZY]~���
�n�5��I�u�|�K&�65��t���R���Ei�y����9��v#:S��@uu�8�S/L6��2>�`��g���2�g>dv�=/�g�]N)�8jhZ��G�]{��Qc�T����[siJs���(�e��(�����t��~z1��aJØD_�d�c�ֻ��� �b�bɣ�<�$�$���c��P��#�<�p]��.�3����9*ݾ����-�)Q�L��4To���b�pls�)������?�;���U�\B���pI�i �H�D"�T@�x�W-C&�|�ʇ����qGAZTs�e�G����&���e6�o�����4-�����RM��`Xu����`���Ǚ��~Q�湚���O��Oiu�yN�m����.d��f�"�����v������g?-�i�냟���i-��k�1?]h�@gY�Eh�7!�/b�/Hp�N���U'W�B�'��Z���3��'��
4ǰ��x2K�Q�H�� 
)mH�Ʉu�bZ�=����RJ��3��n1�;��F��o+�w����N`B����R\D�cGX�~B�$���i��wt�Kc���?�Hr��C:�O��7�F����h)��e��g�G�D�U��({0�[F�7�ׄ���@&�gm��V5}?ۛ�4Xn�����m5�V�*�q�m�������;�hA_Q���f�~���d�zfH�K2׾`�E��_�-x{��7���$�p���1 �b>p-?#p�=�����`Rz���EyX@4�z
Z@�伍p�Z~hQ�밶��Ƕ�����ɀ�:�T��h��d��k�m��)�j>:�[b��n%�fB5+�������c�3%>�%��ӑlmx�� ���E�o�j;(�v����T븂��-�f��@���X�+b����^F�m��lb�?�֯��v�3�6��>.3�=:v�U����- qӒ��l���Yܾ�X�4��� V�<��D��j��X{\�(�~uSW�Nڲ���(��b4�� �hyE?����t3��b�g��X�'��hI{��on�`���i7��`�6��x�HNϠ�D�Ӭ�>j2�^���u��S�{��f��Y��[�a���C��5��`&�˖Kf�CS؀�1�{��cwj*����e`�c�&�՝\�!CY���f��cTTkf���5�{r�8v4P�?Qs��9���]�_`��Eg�xU��gd���sG��n�߰MB�W�6��DY��Y����
���-�����J�-EVU����Eg��{rq��#h0^�Y�1��R�V��3>�4���&�+�r�t��]c	h7-S{y����*p��6��:�d��P^L]IU�ґ�F���S����`��Jeu[xs����ڈ.�g����At���@e���R�}����-Ae�'[%��$n۲ś 
.�8-��3���z�+Ѯm=�2��$�c�N+�@����LK����@!J�I��?�����"!j~%7̀��k$�OI>�����Ba\z�Ȅ��q\Y��`����b�����%���T\�h%ņKc0J�!�(5�H�v���N�M��]�ň��B,5>)a;D�sG"R��Wӿ&_�F'/0�j��0�/�w"^�������R0#*MӈH8����fv_�8��%x@�i1�(IT�1W�YJ��]�%��Z���}O�*�}}��>��� {����ı�j
[�k�@��������<� �~� r�I��mUu��Dt浍�ޠ��Ǐ������SP�0RFv��T�aK���3k�Ԣ�z����Ϻ����Y�Nj��2�V�tڣ���� �T߁@g�-�}"�x�>�T�{