XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��wM<����!�����=���M_�����L�G�ᑸS#��EZ����a!�HT��� ��j�%�L�!���X�MXk���/�D2 �M�M`8�`�/��,-�˯/	��j(>w��{Q���H��
�p�]/�e��
d#���K���AP�`��O�85�A=���X���T���3�bE����cp4�N`���n�2��gU^�xڂe������X���B����$��+�DD6d��{ἆF�]��룤��N��c>Y ��R͠����d��6ݔ�Hy]i~,OK8Q��0��M4}|���@�u��'�vA����`OS�(�^�*<2\���ds(����aq�ʩݨ�|ȏly	�9X��><��@w�謓Kq�q[-�l&��8���������9�;�(����u��M�G��÷i�Q4˲k���*���6'qEe��O,>����p>�k���K�zTS�eN!��� 	t��&�Sz��_9�Nz���/e�U��M�H PK�wQ%����J>t�@ԾN�hv��=j2��&����~���_M�K�]i5��\�'9��J��y7��02h�MA�3�ZN T�jRIGu���v�GQAg`o�V�Δ3ϭ��o���(�T�i����]�}M��mNjo�l%�M�Ȝ[��O�ĺI򂨌K�ʄ!������Е�3�\kl�d��4f۔�m)o(f���3b��JSY�:���R�5M�����b��gg�ɾbA"Y��U2C�;�EB����XlxVHYEB     f6d     6f0I�>��ohq��G �fm���Xa%"=$	3�P!��$�+Ѐf��n�/�~�=�!�WX���X��]a<SfٮM@	�m�&���^�����ƫ�ȲV���)-�b0}�U�Wl���+���L�n�k��L���v=�
�t���i4��x"�l3�1�u4�!�^����SWڃ�Ps=+Y�kT��|�>����/V���nXZ֜�	g{�,����G�&�|ߥ�F�1?����m �v����Z�5~�ɜ�����6 �6�U�ii��k�_��v�_���	75��\��_�]���L�e6c�e�dS�@?s���LQ+��k���"�`F����R�T�M}O���1�dtf5�r8�$ܪ������'�॒Xt�E�^]z ����i$����FP�2eKͮe�z�x����
u��yr��������	���s���d1����#FAm/���򫅗���gy��F��&36��0aR�(N&0�E�K!�8r[z,n�ɖ������w�u�f)ftlp@E��M �Ҥ{�U2|ы������kO��| <:���ћ�u������4\����\���;ђ&
}�F���ڥ��\�E;����?��H�I����\"Å��g��b�L�o�!��\��׉��o��ǇVh��oV��Q���FQ�� �.�b�^��<�t���cV?�
�J��!Q�q��^D5�%@{�5�'��)ߴU���ظ�+T#�ɍ�x#Ϻ�0�r�`���}�زQ�2���e�FG���VJ�q���n[���WC���[���N��Kn�a(C�f�hm#eW��N�H�3��@�2"�8Hݖ�#��-�3|��p���`�Q�J�����o�;^�E9��q.E�C����YO_s3qH�x��>u��+��֎��Ц�[�*�u�^�;�OQ$�(+�l/=K��H��[=�S�A�:�P��`ڪ�;hpH���(�#epf�PE_ble(gP����=��f�@�3�N;�T�[��#B�$�ްި��R���=��R�m]�D�cc}�Ԝ(�E���Z(����,������� �X@S����՛i��Wml{�<��pF*�ljᙖ�em ��i���7���-�X�d����C��RǴ����#*�� ����
�Ko|Z���Ȧv��j&�(���p�wj���9'��L�T�[���ez��֖�(UM���ZH�>�-�k�h����@��O���B�YKe[��G���3����8������=�=}�O�aEI?ݭ7���w�@᷸my��'M���f%���A�b"7���l�Wd�O;���/6��,T����z�.���R��86�f ��2V�l�8KQ�{��Bh4_ʦ�8����Eѝ�&����Cls|� +GF������Q����	�YS��0�fPA��*S�ӝ�������aoc1lqڎ���>���C�te�ߤ��!MJ�'�ņM�K ,H���n��}ҍ����I�6��ɶWD�^#و�y���-�f���=�`��t~�{9�S���@��2P5�	cs���Uh���:� ��u�7���W3Dǿ8���\�KaIr׬�Y�1�;���r�s���Oa7yߵ.�� ҹ.<	�:8  ��杢 
���T�UQσ��K�m��!a����[�����kk9U��i/�#�撏P�[s��&qs�Q�u������ѐ� ������؇��