XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l�aQ3�`cS��i���ڥi��HՏ~W_/Chw�H�W�Ko�@P�a��К�d��ơ2H��!���̽�3��m��/�%����]9&���q�;�Qq�p��ؾ&�k��1,�������7#d�N*wѨ����<&V��=r�B"�g[�Upkcܗ��^Tg\�Ʋ� S���G��;��堕�](,���2~���f1�D�@8�ʏ������L?Q�%����GE`\3������ �y+�}�̧:lr�X�%�e�8N�WN�%E!Pj1�ke�� �[v�O��:|�6�}N0�a3�yҺ���qP��:�Г'B���c��nvHhҺ6դ�k��^&|�[�By�Hנ�w� y���gR)�L���Ɋ��p���*�q�ZmT?9ڝ��@�+}�6�l��[����Q}�o8Z�p����Z���"K�f_��^�ȯ���1m�ٜ~�r�{J>J�U��F��p����$���d�)!0m���CX�ۀuK����RJ	Z~�{���F��0D�l-��e�P1�bH?jPL=Pr_j���S,'���c���;?W��{f TW�L�~�6�WŃ�:J~YW?}g�N����'��q��]���t�2_aca�%����l`���#r��"d��󇀄=>h//J%��.Z6ޱ1H$��/�1�l�FKk��xmv�M3�|C����]���Aֿ?�v#�N�Qz��ܽ���H[bp��1+F�w��ke�a3e�I��'Y��h�XlxVHYEB    a037    1fe0�(-�"����Q�J'^^*^~�IP��B��1��v���m a?1�zw<��#�@� T�\��N�Sά�����_^�z&q �&7g�}����-_��}#���7�����t��R�瑻�3F�JUx���-�"e��>*��V�D���v����%ʿ�O�PR1�hP>v��Q�500�v�J!�ڬ\��;\�������g�	��7���E<������`����;�jF��K���a�7�u�9�
ҷJE�҃ �/U����E{~�Չ$6
�w^.G���C��T=2ioh�OT޾X�b!ZF`��<Y��R��R쉌���Y�4���:x���VN��d:i":�=Q����n�B�{!��4Y�ưk� y�������������q�}�\�FB�:�/lC�d-�.�ke�F>g>j 㥉��[wɇ��Ć����#�H�[&I#E�§$f_�m�N��jZ����#�t39x�n2L�f��"�M���
�l�0�	]�Q����&�eC*��Tk]�ơ#r|��r��Ȧ?^Rv��1$���mAK�~Wx| 
Ux�/�k�>)@������@@����5֡%o붻c���1x�~��~��(a�dwYn퉷����A/9u�<kFr#zE�����ddʀ��U' J�&����p*n�E�l�8�b��:C@I�d.� �H-:;���!�5B_U#������w>��y����yt����X�E&��qi���]q����ϼ�=6c�b1v ��yih��&�Ă�9fO��G��k�DH�Ԩ#�����r��E�u���8;���e���uE����!*{���:�(�vD�d3��q��O�ڕ�1z+A�2#Ԋ�)�|�͍���b��K���t�Ҵ*\�Cp�`���Z!�o�~�gҵa�(�e�����:�I�����
�D�����q88>�]��ao�Mc�bUZ�jt��s�k�.�J�.�ΜY�TⅾM��`����2��9�b-����>�u����SOڪU�\��=��F~ �K(�m%;2l���Bz�o��;���֯	��#��g+����㲽(�V�����kV�r��s;���ӊ<�v%�����\6D]#� %u�]Oͷ�f����-LH�������W��պ��'�[�>�ԙb䎉&��2�j�B��u�C[)^��R��)�6�J}!�!S��m���A?6Oo�hѠ�9�Jq�Mz�Pg�u���wI>�>���H����FW�������u����5j�լ]�0U��J���{��ɏ=ʫ�yaX2�jG0D_̮&9悴�_D\h~=��Fu��o�IaL�q;�Vtq��s��#x���p�Д�Sg��[�OJ�ό��.Ƅ��~����cU���t�̕0+�e.\S$Ʋ�%1ɹ�D]�+�U����/}�5/������	�p��W��lP)�_'A�sx���M�G��^�,c��P�>�c�ٴ*�'�,UUtfv c��F{��,�WX�����b$�^��u�����'�M�N?]��	���s��^ֆ[�j���a�@�m�'��5�
�@:+�Q>��j�<iBY�����{p7��ux�:T���N��h[�a�W�`�Ȳ�-�P�;!��&��
	9�! W4�����u]��a�y�TW�1��iV	���X�#G�D�n����3�X�_�E"� ���k�����e)�F-�ڤE�2��^�m�Q5�q)�qA��G�o7�Nu
�sʥ��3[w�\N���Ln4Υ��E�>�<���%PY��'��EP` ��6�Z۫����!CǯN�q~����nPtk�63������g��v�BRJ�а��j�����ꚩ�KgC<��ǐ��Q���E�Y+��"�In�����ò���/�޺~���B�r�m�s���q$���[,R�O6��mZ��[~H}�Y�z�G�H̵"Gq7��X��̾��a/d�x�(�.� �v�|g�TLs�bWa/w�`�G�<�q����jpL�"V3�<D�>�,����q���%6��+ �2��ȏQ�X ��n�b�����p��o�5�&w+L�/2f�ӑt��3�Y	�g��Y�]��<�Z�M��䥓>���֑M@pY���pm�U"0�+�Y�/0L�#���S�1>� �UF�+�$��BK_������b��P�^��;�U�a�w�.���bN�-@9�b�<xL�6�{#i�U[>F����%$CN&��l�\�=�5�����W �QJ�/6�SQ�s������Gn�s�>�(C���C/��W�1I�y"���:�t�H6����d�q ��q䗇5MX�I�X�I�H��p��s)>Y�S�RR���D�F�m|�S1��O�%]�Qn��l��-�
�/#���B�����q��+9Q��MF?���@G��?��mt.~u���I!\Q ��t���eMl�5�&H����&ܶ�	t'I��=@W�q���l�����^Nj�L��c�74$nj��nl�r1V�9A4S�^�����c	�m���o2!��oAӻ؆�p��aTu�;�)��Y�Rw���g�*�r�'k�D5&��+�νF����5/$.���E��S��*Q-��r�xO��\;�BkE����C�y��9�)��{A�V�d�=g	:c%�kF�~2?2�8��Rg\<�&0�y��_g�q̼�Ah ��#inȢ����&�l�
NEs��N�Z�K܉��p�e����n�8�5\���K�-�޸�^�f�pFGo��rRʑ�K��n
]��� N�u�f���'�18��2�V��n햩�Fqʕ�z�oB���]`��)@���

 ?�.����.����=��_Cם<'�ֺH�5##�,��c��ѓ����Y��Z�����Y��\�L�����F���
��sT5�C�@�]����x���M�. m����?�;{��r+$O�.���$D%��ϓ���7�1�c��
�\�=r��{�8LG��/���8�Up9n�j`5�_ng�i�9��Fh�}	��6��
� �7j�;�3�Xfȁ���B�յv<{:�!�ݪ׳/��0[b�W.��X�d�T)�^�bcB��Y���()�"]��4���/�����t4���h����A�$է����Di~���S��w��D�cZ" ]{uG���4�0L�w���,�]9�aU3�2rcߴ~�Y�n���\��=�̈́��	�8\�:�^%� ځ�A������zp��W+Рl]F/���T��y�����7�N��`��\��¿`��7��5��\��his����L) gV3r��`"T�D���Ǘ��̸M>�����6[E��e��s����-9
�4����v�H/��%%��S+%�a����q���=��l�@_i���Wo�k�d:���i�di��b��s��Z��PRs��=o�S0oD6c�	�ֵ�(�u�(%qVe�/�lB�e�Z��-����.56�
rC`[�)���G�hZ��JS�R;�I��0��� ޱ��֨��N$J�tJǛ�^�A�폜����?��O�I����[�2Rx�x��+E�m��v�p���mE��K�L��^)��T��M�xl!C�B�e���̞O��1�d�:�@���,�^��5w) ��@����E���c�����WhY���
^I����,]u���c����-��,��BT�gT�OxՄ��S��%�0�ϲ�v����� +D�dNn��nf��m���Ycqk���,���)�	T{���I��qT�7�f{�/��ZM�"T� ;�o8��8p���C��GR{�jA�A�zR	��5$�?���x���z��W�$A^
�ML�G[�X^#Ԇ�ӷ^�pf{1�C63�~BB���پ"$=���M�m�B�"��=b5���*+���bwn���i���;�@���yF��r���Җ15�>��ԏH�:\�S�z�@�K"I�NU��C�L]�M~/�x{o��D̰��*����H/��n����A-ǥo����D`h�K���Ue�+��WEC��i�x����>��w㌋텪��.���ur���!���H��R"��{�����|/1�q�q��w(�bgY�]�(#����V 9��R7�i{'�$�8���x͢���Tk\��m9�}�k��6��7�=�]b�8�@�9!���f����v�I���NOɊ�D%�/�֢�'���{�������	���-7��av���N����!������E�g�Yѵ&�C?(f^�Mk����.��n %x��w�/��xo�Lf�w"�:c�a�2��o4�<�]E��:��]�'JĨ�;�\)���#�����3�_r6�-W�q\�9���+��]q�
lZ?�\��k�.��կ��>���Þ�?���!u!�7�Õ�"�fQ�<��l!��?����/N��-�|@��9H�����*!��6�i�bW|T���I��gSS�jM��x�	�c��������`�L�_\JD�ɩLY,8Z��b���&I� ��X�M)�u�@���Nx`3���+Z.sU�b��!$� �Kl=��M���)>�#V)�aR��el|�k�(F.㑋d�gw��Nȝ6R�9������"�XRF^ʘ]}���q��]v섲���t�x�H�N�ۭ[.�7TE�ɒ��ͪR�����q���װ2U�͹�(f=�I+*#��H_�r�/��4P'w<��Qބ�IZKg�����������f#�a;F%��c��>j����z���5��'��r1`Y���<�ӲÐ�RH���/��]�1�121Jql)5ncb3��	ZK.�pg	��^�:	JS�/���qCN7	c&D|����0�Iq�V�C�V:���4��F.����䘨�lp��eu*Ȯ+��դ�#k����Q)�Ug
�j�l� w��-<DM�;�5�.97��`tS�5��E��wf�5������H{D�q��ٚĘ�xh*@�\ay��*��LWJ
������l%5�%�����N�ۦt�΢��>����k�h�bQ����Bڼ��r��a��-%������&�2���$D�������ܧ��)lm�K	^rIb);#6h�����5�-z���q�B��'�i�}+�qt�gaP`;�/�WH{���X;R�ؑ��\i8���M�g"5|�uRl�r�fhe]`��|)P��p1�A9f�J�W�F�9ݿƾhBL�e�l���h~.����A��	_�{����^tx�7s�,�i�HϚ��t��GO�z��abk����X�����X;�����#��km�#��=�	Ma�������&�_3FN'�d���I%l�B�Gk+��<��N#��2�\�-��������n������̩�^�� �ϒSM�~ko��F<`ml���O��-�lQH�M���*�%��FK��xa ��=���TdI���W��/ޤ95����G�R��-'��c사�E�?qb�ЙLi����^�3��>��S�2�tZl�x`TWP+�
�M����+�H�;7��߳�( �Nm�`PX��~�x}#p)!̪7r�yn���q�`5�hT	���Q[�Ԩ��}�Jغ2��0����1�r�w��eI�eksǳE����H�սRP�Oe�bj�u?6�'U�c�g]���ɺrbA��:qS�<zHA��+�]05�4Gz���=���	}ꗀ�b<��aC�H�����+o���By%Hn�ܵ���
��G�-�~���G�MF��W�^`)2��k��).�lK8G��c�XV(��E۫��;��r�6u}���-,�7��^�����H�����ü�OQ6�.�X�ƃO�'�ɽ�/lIZ]��?��%�1_�i�����ɃX�3�}i�P|������5��L�:���B�ʤ�G�1���Xݚ~)%[xm���7�p��1W�E�lb�&!n��
h�
�U�r���W�c���H���Uο�:�|��U���O;�������C.jvVe!���
z�}�C��Ϡ�K� r��<��(<���j�D`���5��C��x�#�)%5�
"�h߈T�Lp|9�?4����x���SY��ӥVP|���m�Qx�|�v���P����ޅ�cZY��*�>\�9{P�Ԛ�K��a�h�ǔ���\��KQ����o��/����:��:&	�|�M������Т��K��}�Ĥ��6�ٴ����EF�����=?���.2�[r����&f�G�\�[nvé��� a)oa-.,�P�q�d�E0q̣�dɑ�)�����A!��#mȔ[^�Wʙdˬ����VM}����"L�2fb����V��L2_ц��2���\$���s�V�Vs�q~�'��P�d�;y��\��W��:�wՇ���/�<��p���G/���5S����-�p���ֆK�
<=��U=a(� E{���̼�Α�+�|r�k��c����D��eΤ�\�.{�`32���MD�K_���-nx��(/�/Ϲ]j�O�ͬ�op3�[blt�Ǿ�����1ɞ$��)#. f��I3v�8h<U�8y��IA�����u;r=��H���
��xk�Q���QF7U�0��g��
7W����Ky{�����M1�M����&��~f��I@���U��d�9{�J���,w�W���X���/�l��|$ˊ������#\
*Tx���P��� ����U�� �����i��ٗFW����:����.괋/v_�j:n�2/*�S22<�kI!>� ���#�p�?�.�dp;|=�6�}�h�GB���ā�K���g�]���|6������w�� �����6�����Kd�?�`�~c���V]������ͤ�^��H�NoV���������g�
6X��RR�{��TJ��'T˭��C�D�'-��b�b`��#���#��C�/P�خ���O���E���B�t�Jtʭ:P�� �B�<Γ�3���׍��{8��lN� eAH���K�ҙ���n)2S�+����7}w�cܒ��@G�[R�
5 f?�_(7]L#+-�d�:_X���ǡy�x�0Z,��R��0[��I:c�&�f���(��	:>x���X?�e\�����<��u��-Zx#�*[B�^:�n��A�~�������5�j!]�G�s�
�����������z��S`�|&;
t��
�7U��)ax�ч9���=�ʶѕx٤��M�(3RO���:���J��֫Z�(ҕV���t�i׳d.=˽lU��=3�Q��^p��bq)KHP������e"�gg�C�uy���O��3/گ�jng,J�2�C+w�5�6������SL��`p����ְJ�����:�8F�v�+y6�!������G��E��Z� @n!,�豔:�MBn� ���I�Հ�7|m�<ί�+Z�����I�$�ml�2# ��sf�Kn��F���_��Hqc����b�"�*����x�b��Z$����}N�fO��5 X��J<��#-݉�f�]��(�M�A&���U�=;�Z�O��wi�6t(�	h?����ԇ�u/�f�ڣV&��x���R�
��v��G� ���ϻK���mȞJ�9RZ�в�������&���-=��d�W)}Os�:�H�L2�OF�-��DCx��I;Q��Y�92�!фK$��j������|�'�}���r ����M�a��%jq՚o-��߱���j��;��f��m��h�ꩊR��FO����^��7�܀�u��b�q��8B'��K��ve�8�A�hT�.� v���w��m�ET����T3�9����m���DЧe�	�;�|�E��#�=7�|n�}]��<3d��������o���r�����1��`S���W&&_qK���+'�2a�\��,K�-u�����6�>�nvl�!��?��(��[�&��8MQ�&@�íg�����^���!�G�r &Fc6u��<���3�