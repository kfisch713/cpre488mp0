XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����R�ۏ���$I�"h?�K�A|��}~��^ԒU5��߮+�qo����E���'�/�^���� Z҂��ܘ�=���C�Aw }o�����Sб��S��\�U��'����))혬M�M�U3�<�<*�|41h:�x�?H\�!='?z�P���m�-Z`=a���Y���)�Ow�~�`:�cL>5�7ۃ�(�\~9�J��1q����v��𭬫�M�L%��>½��^(�`령	�]���T9}MK|,�*s���G2��Րs�e�.��߁9.]0��p�i���|M�����c�E��2������Q7*#�]�G�m���2e�9q���^&���M�%��_�Z@SF��FG��҂������'�[�3x��T��Ȑ#@.�}���4ơkaj�W)�� ���b𔅨s�2��}9��df������A�L]ګ��k�r{���R!�I�+M���j�[�������
Sw�]��i�C^�$ހ��J��F&���m�9�B�ހ���*�gw������Ѣ�;��(w�]J�˔�Ʋ i�ɕ��$��݃�N�qa����n}�d%�n�ʗ�O��̳��,S�����Ă�f�K����s��.���Б�C+��U�����=�޴��k�ٕ`Tk��w�<x��]����[s��| �E�\R|�������n:=i���|�;�TJ�}�S�ݨNAF* L|����Gb`g�`���OL��X��|�{y,V��B����XlxVHYEB    42ae    1110|����'�ۀ�����v�f����fG؊�J=ܢK�C)nvx�ek�*+r��.O!,�<�l����.342���L.�1n?	;+������͑<G��Ñ{Z�y�uo�-_\��	���ohT>��~�4��Yۢ�؃���IE�<H��)�A=7ZJTcŮ"r�����}�ֽ��7����e"�Ip�M��J+ں�X#d�mP/�SY��EDc1���b��`O9V�l�<(2��-�Ű��?�B�[��/����5dL��.#S��5���%V|�U��\+{��j)��LO��#QQn�pWM�*��k?Ι�{z��ߢ�U�7g���o��L0��>jE�πx+xv��ќ��7��knM=���#�a���i���b)㩗nȱ@
p��P] }���(��Ay�1��/�z)uZ��7�h![�y�SDe4��6��m/a�덣��/O��Ŵ"P�"�K�>$��N\M�n��v_��������ӡa��	џy�Lp��r\��Eq�I@�a؇y�(�x��bG��z}�gq��K���n繮�Kƪ����{ٗ; �R蘿M`�UH�,P�]�J�:�(��/+[�nM�`��d�NU�qՅ�Ŝ�%��^ >�b�H�O28���+�8�cO�寊T���P��|�Kh�.�&�.�]hN�pI��Tt��s���[s�CV���R�۞��#�#���N����W�AAqMg����W�; ��ʠ��⺗[Y�3��`+�8�C�$���\��[�u�����n6 �i�`l�п}R}��v��l( ��k.�@:3r���\������~V�_H�*��$��n��<���A9�g>�4-��7���)�8�R1ػ�؛Y��u~R?����3�i�����ۙ��:��C����_�$Keb��یY�	�����|yA"�M!�2��#$i�ԣ�:��e����ЪY��G��A5�aQ��ҠbC�:�Q��rXD�+�
hf���;��L4$�X?��20���J@d �,f��à����g�e�&��S�~��?Fn��d@@�t�+�~cϓ��$�	G�q��@e���h!h��/��'p�H!�5�LD�Fk�W��>,'�ik��u\�W��*)����+ڙY�	;jW�9�7`�D8���Pa��-�C��X��*{(q��	���g���xkt��{_?�>#^�l��j}�ID�tCVP|_T|(�`B�� �F3�8��Q��?����@��`)��2�^�����o#zM-��@�ǎ�!�t��'�Cy��kY�K���g��� �r��=R\B
~����`�.�J�nd�SL��宝2�\���U`�$y�_��e�.m���2;�"�u��������b(�ۅ�T��!�Y $kԔ��?$i�#RA�	�)#�{����|�g+�.���� ��v����Dc���B"½%�-�/�����<�-�}	U�e ����D��m�Xȕ!��0�;Tf���8�x�"~3fEn��Z�7]������8��41�#�XדP+m)�z����C�� ���6$XWuҵ��v�nJ�T���Y� g��
��Iy�M)ߏ��N��>��N6'B�X8 ��~)�)gb2���c�kU:<I�Ǡ��ӝM��F�N��ޣb����%QBB��lOoM��������s}Au���o�o�YǏ��[FR�K��>��0�}����֒�Ґӑ����(�x��%M���E���7�.K���Gw�I��c���E?}�z��4n�H@W�m�ߺ�	V��yߒ�o��)���� Z������:Z:i�-D���n�S�M�5�D�N�MxŌ��̵V ����p@��0a�CcQ�� 6��GЫ���q����]_�Lrѹ��a����X�Ȧ��.S�һ�%�]�T��.r3�G�y{^!���3�ӧ��hR����$�lhrAېVg�+&`'>�=�v�=�)K��c�kE��Q^�qv_6�ǃ .��������!�)	���[}��+0��Y�2^	�1,��u⣌ق<�s7"���W���0�������!��bu��{H�e� .��~P:��EF�H�@��)�T�@�&.��E�
�%�����t��9��zX�^�r�R(���.�Ř�Kc1�����c��@><�.d&��5�(�[G�-!z���$=����'�>�$3��a���9���*�/4)\O�!ȼ6S�~�ބ�Yk�o�#2����1�.d�q�I�aȽqX���*���_�G�]|D�@il�(��aTi�N~hTz�WhX�.#��ZZx�;x��PBLё�Z�0=OY�����r`/�-�4r$|��#gEJ����Hz{�+�\u|�n����[���\}H,e�`$d.��I	��f$�C`ɪ�ޠ��A�:�&-���I$��.���d;8y	��1z�z"���Z�U�H��-�@{�+k�b�lIg��������kD�p��i��2 �;�7�ƙ�؜��9k�	-MK:�Y���E~�`�EQ儽PF��2{���fK��]~�N��eO0C�8����d(�>�PG�Vd�t�.��rިU�7��s���$�Qy�~R�ts��Gx��T@�:*����a�\s,�c�	��	kqT�ܞ�i�7\E����F�:7��&iT�v��!x�_mZ=4� &p����t��Ԩo8�*��@36'�i$���5���a��r��zy~QR�q�{�0������>�T�o6�P	�e�9%��mpF��:	��w�ԻM������ɉ+k+��!�z�1�:��޷����v�gէ���;�p��)XY���@.�wl~��KhY�M)ALL~��Zǔ�+yO�Ɯ�!%Z: �qK3ทg����.�~����eޖ�:ʳ�/}L�jtLCjn+�i�F��²�%QP� �5�S�-��j�99�h���d�n<�2�k�>y��Wk�Ti|`�J]om_��O����������̌�m�n�����T[�j�S׽TM�T��vy]9���x�ڸX��X���c#{p�v(��O�Q�R�Gc��eO��Qp)��f~?E�;#l�	HΨ�?rUZ��Ƹ��̓v���/����V�1����K�˟�"zo��>/�˖�r./�F��ņ�KB��NT�����"���r9�N3�)��]j*s'鏡�^�1;ù��[�����׳
r�ju���T��v��к�0���Iq�^� 3S���sI�~�e_O�x��5Z�N}�2��>��	F�k�������o�������8�MA�����j��ڋ�a��o���-���o��ה�#�!���F�K=���h���h����~��]��p�,���w%�I1�_G��q�	y�����.a��;i�w�f��y>��n���6�X��4�ɴ�����p�r4��}�H�:������n]�Z+~�p!�K��c��_���Lkϙm�9ڬp�j )�':s��ա�꾒H_@�4-���x'%t���� h���
Z�� {5��جJ����O3�fpn��H	S�nf"���%p�uG]��[d�{����r�e]wy��
��A�q���H��t+���s����wrr�
�����Q��ud�)����5E�s�9�EkU�� �Zׁ���>�1�)T��B��c�x��ޘ�����B&��&���Y+��+i�1%s��-��'��g�K	����܋d�k��@��G� �!��6�:���Q�ɻ��Ϻ�Ć��K��ۺ��yo��s̽K%�Q9���K�1~=8�M�#+ϱ��=y�_}X��5L:Ćk����p���#����v8,�3@���ڛf��V����z�p�C��*�jK�Y���9��^r�����l�O��ئg���g%��M�8���[8��2����<�:W��!�����"���ɘQ�3q��Fv���KuG���nxg]fp�Ѻ��KA㺟b$�;Դ
Ʃ�����,����eHE�-�cI9[�9�̭�ߓ�a�(�9��/���i@���p��Z4�n���u����&�ҹDW���@	������K?�*�98�i�\Δ�֍_�'�"70���2uM~U��W�]�<trJ;�	��4pߊ�B+� �����k(��[z���컐SU�}�i(�:Y��(M�g#�I�k������ �����A=D��v�^��L{��u�_�UA�#ȹ҆���)��< ��L���cz��M�}J���	�