XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����[�\�:.P�n�V/��k������e��c(�=A�5�aq��L��A�{��Ђh���z��%���m$N|��{(~��+��ć�ک�F֝+�;�5�:PF[�7�6�nl���t�󛅀�+(��"ֺC��������n�Y�Z�5�RV%yÃ/��
&�=Ѧ�5�a�Z0h��,.	�@��X�`��]�-@����N�L1�-q+�d��Sv���R��`��h0�ƛ0�JA�x��6��lSO`��er��v�B��`/����x�md�3$V���GuPl˨�����"�U�;�/��Va[�=��s6Y�Ѝ�?'�Oʊ�I	�y��lB��@Z*_ �Of� P}�X/�S*�F��]�,`!�Ycv2����n�Od��g�d��r"-�}���7!|0� �p!�#3/(��ij�)�%Q4�Q-�X��������A����?��f�j��7k�#eM�Eo/��� ˾Ś
�7t)�N内'��=6�����.P���)q|r�2(9E�>��?T��H��We1��NH�Ƀ�߷-�"�cո��v�d�g����g8MzĄX��O�ue���_2G���`:w�+�!)�Rʠ���~���ʄ :KN�-K���Ʌ�/�r�xԂ�ө�u,���t��ȣ�e:�Ce�qpv��?8�# ����-p��"�E�L�5��Ň]a���_�4����({�"���=:����g5ZO+�SV�����Z��E�.v	� ��g]�FlXlxVHYEB    3fdc    1160,�q����Ӣz�2l�s�PL/*�g�:����G�Q��+w1��|G���,&I�,�"�.��Rj&�	����v$�v�6z[��&7�U�Y����|);8�;��a���x	��ى$^;�R�両G}tg{��%q���������W��[���XJ���,���a�:�~�Rv��.���'�k�j�6����ݹ��5�l��/cd�pV�{��ka�R~^���o$�E*ϴp��*J _0� ��*`ӾS�d7�w7�IP ���� �}��u���F;#X?N��?!J{yV0#�;�X�/H���u n-ȕɣ���4��@�n��
�q?�
��&N� q�]}���<�MZpQU����؇�7���"E{�,#�иDv<��gNf���u�z� R���V-XkA���Og�T��8��qV(��<!.l�C�z�o��rX��z��!��/|/��g!�#-��v	��Y�J���ӷ��D�[�.#E�>�-1�3��sr�]�j-Qbm�x!����ڜ��H�.�&�ķ� ��Y'!j�P�M������䴸�˭�([[z�fq�7v:������Xz�(�PU�%:����>�Y�F��S��]�YZ�n%��<�#,�`���&&RtX4���ܿ����+�L�X�%�~����p@q�>|Ƃ;�`�|x���qf������`��T��_n�"�mU�
��W �E��U�-��Թ+y8 �'�i5��S?�����W�.�kB	QmÌD������}��83G�g5��� �t�G�}[yqFV+Z/ݲ��Ԑ8�NZ�(�@������+��6;����[⠼
,z������|��A!|�H�3^�"�(lͺ�~��QMN̾w�w���7h�t�7ă/��Z2�j�,R�i�O\v�d�QO�,�1�[}���V  �.���S��Q���=	°��.��V��1�;K/L�f5(�>9M��-{>3�P�u�`�	����3�0�Qr��DF]���p�ݒ
t��2��gx�S?(~l�$|s���ɩ��K�ϸ����I�z{�g�q�,|��	���Q`P!�u���,���IF�����(�d��Y'��g�ߋ�#�A�y�i����I"�'h���k�C�Y��wM��\R���c ��QM��Uܥ�~�/~�q�e�l�J*��$gq��e[k_�>\[�K���V�C�Cz�J�7{3t�@	Z/��pE��帇J�t_�,+��u��$�Ֆอ�2�'k�tl������d��u�~�~��t�_��d =s��X�߽�p�h�lā�Ze��Li��Q�z -#,������')���Mdb��k?�Tz;b%(�Y��A'ʟ�������{���3h_ѻ�7Xk+��;�A�H��Zӯ�!�Y>vo�eC6�F�t����B��qTS= f'�Uc~Br��Q��Zo\���2~��ėԮ��o����" Jf�eEU����8۰.xW
�en��*�D���q'���u?\�+߱e�^5��xDJ�6Ԭ��&�n�-��s����	K���@��Y ���Tvv	�Y�kњׅX��1mo��EW�;��"宩���Cs�����J'y�$oz��uzn[�E�=f�#xP�Z%�ept9���
��۬�g�̖��;H29c�i��d(.�����K�=��i���ў&9��%4��b|Uhp쇔@�'��|���֯<��֡��Z@���Y�G8t�iI=�d����1v�:�����ٴTC��E�)):4]~��|�uA�C��ʶ��z�0���� �r��_Q��-�r֪8TO�o���C"���ł�=B�58,��Ǝ��ruH�]b��J	5��T�~�Dl�ئ[��j=�Z& ��.ʳi����3B�Y)�t_0�8���=�蕑��v˦즃�	��䣷�"1�u�p��v�~���{��<���E%s��>�2=+x�6�#�6��H�R�XHՕ�_�J�>O���c��|��������i�Ȋz���$^C��*�(��-�s�|Լh]k{���Lʝ�������a�E2t�[6�~�[�~��䃡���M����^�Z�kF�|��1qL �ԓ���.��Y	�0��9�2�H{���F�&C�3�^�m6ɿ�Y�Cx��'��5�]z�����n��&X2m��_�7�9YZ$Q?�?fE���􈀸�.5�� �d�(glV�?4֦fݱ������Q.y9D�^<}��H�R����[���f @h�f9�6��.ǋ�)�^:��S@-j��9����e���<��O&d<Ly�B��{����OX�����l>����ui�6���7�[�����։�w�?���jz�+�x��*���lp?�����e<��k ���������-&��GO��x�;!�B`��M.��+���\��hc:��{LC��c�@���hk	��
�����x���f�L����8}�uZ©�z��d���%;��X�%����o3��(���kg�<k:���0X���u�e�6UO�	"Hԡ�RP{p�?��a��F*����AG�7�O*]ǜ��G�u�N����C7�:��}�JfR"ø�wD.�j�@�q���`svC��k���%J*ڌ�6��RZ�/WHT���;k���Sp慳�K���QB1��\g?n�YA/}<M�1G��;�x�B��`z�b�V��4�)�yl%
����$e=�i��f�n�Xs�Qq�U�\��}�!%�D,��yVN\0:��$�����r���9��oD'��Nhs��o34�����-H�||�-Q �B�Ů	"�H�A������l pE���g�3&$�(4n�1<'�nY6���m�>��-��q����D�+������ ���\�֑�Y��K&E��[�|ƕ�@.�sD@�`�D�� �t;�_�$3_~w��g(o��C�����΀Z�šH��!�%Þw���τ�۹�W+�
,�h��	�����ۇ�A�=��6j/X���a�|ٺ�N8�}ctZ'1mG'E0?�f0�M�Ძ
,ˆ�'�dw>�dt����{�ܪ�H�m���>؂�j�\��"�0T�`Y��ȭly�8�|n3 	U���\DB,TM�����k
�3"IT����&p�t�Iz ��`"}[�_m��}���ؐ�7�K��g܂1ХU9�6E��'Ņ���!�E��k������ݡ�+���ja
n�k�4����j��ƽ���G<����� ��X��W.G����W���4^��9��oNL5z�$����`��dF�8T;2u4�%�Uvt#@�z�⒦���I�n�.�of����c$K�[<�ۛ(�����߄��\Vw��lդ������܌�Ҭ�ү��Ɵ�m�]zARIzD�?����N�L�^,���sz{\�b��.���u�B9�aس^Q�}�CF�^Lper?�����ux�1��#U4�Ҷmʥ���[����p�=���aZ?��8�D�M��}�U�r�͏?7�c���-i�5L!����aO�R����.z�/���.qTDcC��/N�����"�Jz����P�@a&�0�wOE��L�P;�`��'�(#i������~AbV�ЧY�Ϋ>jZK��Ibiy�2SleZ�Y�y?�L�l��tT�^�)U�7�� �2���I�,${r�Ќ)��[� !ס�c��/g,�6��3�x

��<3S�p�z�6Y���%�t��/���������ب}ZXbu���
�I�-�&	�t��;��e���GQ����&�>�9���x�T:Ck!R���ĹPN(e�p�c���1�Or��z��̻R0x�,�L���QA���@j�S��h�&ފΧ|c� A�yaEnԐ�z��Xe�_h����=�[G�,�v
{>�4A�����n[V�(���+�s�Ӊ]�5�S�X]�8�տ{�yM2v�R�GŠ `r�@Cb~ff�������Ic3t��hQ�{��c�m|����)�kK����$du3���hG����YK��)��b�vJ�U�[u����2����I��^<
y��X5d���K��T�s�[\�Ap ��qR��ߙ�ݔ��5��]�
���ԓ����V����t �觵@�"���z7�9Ym,Ȫ�x��V�Be�A�N[�,�ٔ�~���U���^����Uy>1�VC8Rn��bX<�c4���/�Z����}��� �J��ry���*�@�7��W�-nkɚ�YMc�W��D�_�a���-JƋ�vA������o����&3�M$�Ĉ�?�'.=��G[��k�
�u�y�p��B�q/�k��yed�j/r�A\�T[<��ACS� 0�G��*