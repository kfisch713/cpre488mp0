XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ۃN��č+��1�})e�2U=BN(� �q�����8p�s�\ⷮ�KMF��׮ߟ�歏�u�D�� 9Qh��Ⱦ�D>�:�h?D*��\ ��+bkT�<��{d:�Ê��+�v�ܑ�G�9=��ܾ5q7�Y�f�*o{�sK�����68WK�
܌ö+p@�	Y��6*/�$���A�~���;u��z�/Ix���6B�6l]�&S�xP���b�z�![������'�'�įUS��������7��3�r��˻�˶��T4���
l̎�r�����]���tb���g���f]m�qݢ��K���ᱬi����WW]�f�d'L�H͸����a�Z��Q�:�I����Y�p|��1*V$HFl1g�"�Pj�8��G�^���R+A��,��u�|�KH�1 �+T���ēI�8n� �{N#�B��O�pH�{������� �^vN����eR�]���Sx� y ��c�g<`�z�x�A��*����fᡣ
��8��uz�Q)�H�y���w�u��>G�AEK��胋�+,HR��˔g�%4�Wd#`�_.�l+��,sE����f��>�LX�L�O�c�H�)�ŀw{����xws����9�2
���	��M�k�<\79Ҩ��>@�C�{���6�6��흘����1�5#��;�|W�h��S�_(Ѩ���r�8�LY\��e���ϻ�G�)�
_XlxVHYEB    fa00    2040R���_Z{� �:OI�K"g$!a�-���K2��J
ܷ�Gxܞ���W�F[��_�0	���on��,Mb�#�x�&"̨��e�Y]�^C�L���b#RW�X-��h+ hw&΀��e������=��:2��M�`F�����%^�L��dP�����8`�l�Kr %{����"AӨHx5U>̓�̷�zW�(�HF��k�D���T�:���*�6���|:�/ȴ"�`�V;�)�0Uy��օ��O��f�q@���*����麤nC8U�rǲj����nK,WY�4ذ9��z�����c�R�$С�l�R��z�u�G�F���$285~�_�S�%�=��q��n@n�\C"�Fh8}�����A P���FL�,5L�S�%�q���޲>�����\��L똌���+U2�j,!��=�ƍ]���7�.�އ���D\,�J��j� �����j,bn�]����	����D�E�a{7i??a�sd�@s/ᓻ���6�Ⱦ�-�>S 3�s���n
��P��uf������<���I~�*�JP9R���!���3:�F�$ĺ�2�U��|J�]��ڥوϤ`�-;_�.��l��9z�����6Z��T��rQA���#Fݑ3X���n|5��Ff9G�9J���
=]��04v���s�$�������°X��s�Eryu.�%��r�]<DѩҔ�/�8��`	M1(^#]N�J���oP(���`�V��g7F:q���R`^2��P]��1g�lV��t�>����(�K~l��*���qn����tR���mF�'H��I@p|^��\�ȶ�<� -��t�S�#,��ɗʾ�"$e������@AdRؔ]���v���%&7{�leݾ�*n����C�����N�"<6R������?b�6҄����jhז�ug�����'5d�w>��HK����]�X���\������.�����Kh��;ۺ5�8[��:9QK���+�4�(>a�V��R�P���H6�4G?w"�߂Ųc�1vn�[T�9b$`�i���W���p j-�?aHKH잖�Ӏ�����U��s��	�pL����#�D�|�N��B�XH���������"�L��E;5c���eOb�WXUP��B���UR�H�T,��y�᜛�X{���3��@�}����ZB���s�Δ����S�9?C/��@xY������͛ڜh���s�|��Z�ߦ_��Ѵ��`�#�ɛ�:���|���HA��ፎ���,�E
�
����g+��H�����cUtqut���>>T�Fڑ@��<�p���\	�t!N*���µ�_����0YN[O��"�����=}Q�Ͽ��b�<}9E���s���4��p��Sn��x[ޫ��1���ᡏ�E�r�����4#���Ԉ���Jx=��=X�#�����2�0ӕ�!4'�����\|t���%9�����E����b�����+���g��E�<MA��T)Y��Wt]!��P�~����[,��'Z��;�Pa�QzP?�zB	o���z׫�-��m,K$��ƍ�+�0���T�#�Ob�6/Ҋo��e�D��Aq��$�,�8o�@�"���h�J����o%m���cF?����ȩ29)�!M%�t��f�aA��(3�"&1�]��v~�v�l���
^�F9��^	��6u�1�>�7������F�*?�M<�f�W�4�2���������8~�A~����~P���!��08�
o��c��D|�f��Y�Q�Emc?����{�J��)&m�2��*n�(��x���j�2��!�"��Wdn�x�_�~�g�=��"��6�F`3�R�Y��4�&�ڤ���Ϲ%���Ԋ��)��/��?-�Pm�8���CT���4a^j��y����o����ui����HZv_�@�����;Z�����
 7<��:�?�ݕX��D�^6G�p2�;'�'4��G�cS �na���|��r�m�@uw������5G'�^��EX%2�8f��Ǣ7K�5�q��ãK���U���~dgj�]4M9��&�L�ݞw���^�,�a����)��-n�HEip�7�F����1E�̝N�U�Vl>��2�TxGj%^�:<,��N����Kz���崻V�p|����	�t_���=�W|Iδ=��'��|z�@<�0�K�O�,$hA��?��?�����u֍�jͷk�7T�D��&���K��K����a?�Cז#hӣ�g�?���H�}9g�@.�cwL�6|�S3��Fc�������:\R�w6�Dn�{8amV(�H�4ح!%ٯ���-92�^�p��6�&�Em��Gچ��������NI3J�>ޘ�s���ܭ���?���w�+����Q��`,�Uȅ1���L�N���8�7��ˢB"7���6��g0"N�7��mv��^}X����^�m���an�'��:s�F|d$$U:�Ғ"�j�J��*���~)_k����i$}�`\�o,�vk�s�\7�.�/�q$��K���,k��"i�a�×�2����5����oT�!gZ��P�xN*��,�H��{)�-c��dATfj��YL.���@��ГK��E`=�*L$�ţ���Qs�	��k�o�������hc�@^��Q'�q�eAxsc�a�f�����k�=�0;�����0Й;_N�ڹ���[^S�k�(I&7Ig�J�@s2�nz��q/t.)&3��X���4�w�+��v-A{P��-��:�|���6q����ɜ����]��3�"���-D�/1p��"(��$d����ͦ�O�sO�L�a�:Q��i]�<4�
o�I����	3t�[f6eɖ��.]�㉸�=0�7LΜ�����-6����U��[��,�Np��B���&C+˪�]��i*I�P*��D���[�  }-N�UH��jK�ŀ<�/iR��A��ȸǮZO�DN1�b��sI���?�FK ]1��G�yTHt̵&�+�)��v��5Τ�i�V����76x�����US���fPq#L��O*�;�mYB��''0t=��B�G��#%�$��]�#��~v��+s��U����PdIs�Ġ�k�	�xG��D"�4I��,B�̝W��E!>)fc4S��W�\��Ph�}ojڼ y�8@�׃�{yͲ%>���P ���������S�S�������PN
����e��x�����&�1iQ��ֺ7�-�u�����S���L2Ϝ%O�
�O��e�*XX��{�o���I�$�KG˼�)\�z��H���'�b'k�%�g���>�CD��΍cۙf�渮0�H"�T�R�^���7�"!b��K��>��ۮ����װ�s�e'����rN	AZI�Ͱ{��3�ǖ�'�D �����P�!(t 0��uP��3T����E���05�xsm�v�\_�IB�w߂sgT��z�*t(�P��Lw�d�L�����X���T)ZԶ���`�x�	�ob�,}g�~��<��O!�f�ji��)�X�_z���7i���#�j�GG(V"R-�\�Wq��k�?�~��id��9�y�>��B�9���*�W]��ˋCs������
�ÑP�_��h����~�K�q*�RW���l�xFɐ��'q�A�v�qn@˥>7���Og��O}�1���DT�"�)��Jy��(�0vq�XI~�Ut��m-qņ��<5~͍��uu(�(�Jp\M�N�������N�Mt�E���( 
���a�>s�H�țĎ��.�y&���i� WX�����E��g⾵` :-J�~���H �I�g�(x�%eP�y�!W[�=-�u�D�'������r1$2N!Qg G�X��HxYeW����.�h��D�vJ:���]j������	���i�p~��KY�ܛ�p{W̪˨[��dd�������r���e�rW��˭��ۮ@�I=��L��a?{U
il���~�(�@Is˲�# _S���a��A���z�`C�h`���z]�ևR�Nc��ھ���ν��K�2�n�S�gHM��ʴ��k �+��־	���z0=���a�ҽq���e��<C��6�za6�U�2ѱN}�(�ꖜ)-|1��ja�zP_,i�u�l�i�߁�?<�_��v>p����j�KtA�fR�C�t��X�!1�a���T,�-�N�&��J�I�����|٪ �q��	Ȼi�W��Q�b��S�!=Q�1
×����b��P������S�j�����w}��M#rَ4x�����ٞ�M2!:08G��\]�`_�����_�]u��\ֆ��*0�3,��>�Em�8�>_��z3҈A����JG{�l�z",L_�|?�܁�i!-6����s��ٷ�O����y#{��հ�w{QN7�ᦕ��O�Z�Z��ϕ:_0�M����
���(*��v�Y�w2d�@�E�[@��,ѣ/��B@ZC�=�:���2�ex�'g�}[p\�R��j���i�+IB��/]z��h��u��'�mX�}r��rKv�uv�6u�����,3�Y �/?�k�y�O|�/"zu`?�he�P�@�<�p��OK�W�v��$s\����ҥ�M�d������2'���CO@��Bl�*��/'��9����M<�7�v��֛ь4]dd����W7�R���U��XV�b��T��H���Ǐ8��7Yl���i+-x�2�?M�#�-�]�i��(�M4�ޕ��e@��u�AӅ����6��m�Ӏ��������E��7��=_���'(�+�hB�I�F�ƳV �k+���Dܢ��8�ɢ4ՠ	�&�t�_վ�ΚÁ�38Xk��Zq�(�Ҹe��S0qz���}�i~��<w��㱘��/����t���a죠�VЕ�����꽚6�%�O�V�h1./�Ff1k���6��.�*x����*�����C0Ƿ���-�NDӗ�����R51��գ�*#!'6֋��D2Ll�v/í!�^��+�M�=)�05���d�~q�I���r,�4Ik��nX��ס�M�r��>�:,��L�I�z�������}/�ӭ�Y:�8'Y�;�k0hߓ��ǂ`��S�h����4����hT��(=���H�X\�8��%�6�|a1m`i�}��:\�:s�y���$l�@\Q����Wt*I�\~E��tq�'Μ�=y4W
���	�'l{�	I�* �:t�J	
s��|��1����?�����zT������g�l�;F�V%�LJo�ސ#Ϗ��E]�d��Q�3��,*��%;��ÊfIJ�����5�Ua�$��hb
�d��^�j��t)�:�#�*d�i���Amr6�1�HL�'��#5�����@:�<jF�b��aG|��Z��V�n�y)ؕߨ��29Z{N������qTs�jS�����Uڗ0�n>`���TT����$v4*�Lk�����e�Ӥ k��IkŸ������h�U`U9���u?^��~��ؿ,����R�K�BP��~W��F��1W��-���� �~mL!�0j�ªO������bw��3 6�V�=Jc�!um�N�ؓ3���"�߀laY
�,��-.�-H:n/��O���U�C^qޏU�!���e�~�@=ͨj�R#�q�[�k��$��d��H6�2�Z��� ��I{B�`�8q?����v0���@d�y� vbR��I{`܌YrT�ƽx¢H��C���X��!���c+g�@�0"\poo"�"��~L_��>��<d�,�0N��1��Gϩ!~�WCú��<���9�٨q�`?Y�j ]"<�?}����]D{��id�I;U(ªkk�3-��h�l��Mn��n
 �4��V(�~�i��tM@DIm,.��x��b�U�'4d>���{5d�&$��P�A����x!aP��O��枽c7:d�5����G�ӛ�&>����&�W��tg�cx����$���?�Zzxg������|��� �HF���'�t�_fL,���W���Ֆ���Zͷ��p�-�9xw�<����d�d�%�\<�ڍ���,�p]��������l�O�䋘����(T (�����!�X�tF}��x��\2�X�;b�qŤRM?(�gNNUY{�L�i��G�<>����W#�U#Hf���o�u5�rj�.��&�Ǉ��p�6������O����"�R �U�^�A�����",@��G��I̱��o�5�A��o�Y��,�Z���#^�2T���X�p��߀����}�n?���Q��� �_�	�N��XS��}����f��pqW����F�[[�Ŵ.��k}F�	��#�ww�I+2�O��]%?f9]����k��΃&[�}�к�J����rrfq��Z�"�&�.�ygF� P��D��e`����dN��{��ͪ'���ca�6;}ұǼa��^���IF7bn�r�Y����b�N�M˚5a-�p�����f:\R�N�N�
(XB�x���.�gxm��¢�ާ�"�_��+?���]p��L��N�F5�;Q�>H�p3�"�K��� �|�ݓG��a��lfX��EZ�Bh�8��R�����7��W����i�=uq��O��&�y���h�Q���)>F#�z����*��A);���Գ+p�����>|�k�QU�pP�	���v�����"91E��u5�Y3@�)g�����^0��n"�p��.�B����T����"S�q�tc�4 �(H�8f�U��g���Kq ��|	˞�-<��2��2~<���w&=�yJ��?鸽�b}���Ɛ8�˭�<<��Z��9D������{M#�`	�u�0�O�C��\V(�k	� |*���p��j˛/��<�h��]�ÄE���,��y���xQ�}{���n�ksv\C�`�a(cU�A�|D02�
�����̸*2V����J�6ۥ�(E�}nJNn���� ��/���_��9���P�1�F�Y���H	��kB��-4�ް��o,����s����O��ɛ���kɣ �b[�e|wKޗ���y�c��e�킹8�}�P!���	g\���.{�B{�X��/A�-k�F�#obR�EH�K����BQӏ���5vn�jX�4: 5�q�A���N����[$�wT-1��5]�K�I	�2;�뎾?X�6cγ4�VѸ��I�E�h��{o�9*K��	�r���3(��2h���@�^�$��1�e+@M�{�c���"�� �}�+��gF��(�#B{�t��Њ �´��JA�pxteVd��|m� �O3Îe��Ϲ�\]e ����Wv��::�����p��]F&1�������+��P���l$��O_���ff�>����? �6t�d��L�?������Z�� DR�k��l��<zZ\:^��1[*�ey
�UJza��Zay؟�0?lʧs�cd]�Ӽ���S�^
:v��S��ʩr$���I�_/u�ڰ-,�}�+U�YgF��[���7%�"@�ϕ
��V����i�uu��~I�^��
35�9L��J�i�~�y����w�DlW"\� �t�~S_����&B��tID�׉cu�Y�A���ǯ隷����j���?<��A��<�Z�uϑ�5���'ODF�8�K��p��;�����*�{���K�5��;vy��7�v�i�r!��^��z�ea�R��k`Y<f|7��%�g[�]��/�4 �=��k]�ݵZ5�A�*L���QS�@����-�h� ����/O��Hl�o��m �}N���l���1X��&��epQ��<�$ҶD�22,�X�؆�7o?�{:5�f�}�E��}m�E#R=L�,>��)Ẹa�穘~�n��G�[r��Ʊp�^2��=�!�/�;��e�`����t�َ��./�x}���r��r����0c���i�]����w��������-����MMkQt��+��!w���K���S@�*�i�Q�k *ŧ|W�^�1Ɯ��h�h>��a"����1�XlxVHYEB    4f62     b506����N�WA���"�Z���tܭcp� -����]\z9v�#����(�������� �*T��M��� `�1�NBr�M�Ф �9r��z%�[)�,( M�,�b��9@R�C+u��&	f�Ç�����0H���cSwX'���\GB������v2�8@$x�|��'����\9~GXF�� ��x��g\H�e������$��q��Ce���3�x�3M�au��Y�ô��ĆfKr�fӖ��ʝ\�~��z�[�"<���1!��d%������:�B�R���,ѥ�,���R�[=Ghg��p�L�뾑����㸔��u�W�n��?�I����h���g�3YB������j�s�l����$I�'Ճ�c�>��G �&B�Cfz��껥u#������1������c"o�ֈ2��ݙ���79�ݐ�|!�T��[Iʸ�u'���z����[������-� �Q����Y&=d��Zc�^+k�;ԡ����ևFDu�k}E�f#Q�0�$k�_A%��E�O��}͓�"�T���D�@�- i�~��wLo+�g6�W��<�k�|�$;c����3���d�&5BW	�!�BIj蠵��
$�af��注��&���{��H	&X.�w���~Y��n��7rD�3"�;�B���d�?�8�h�&��3��!�Š���8����}̜m� ��
#�5��*�<]/|pGZ�����[�H��5� ���3HEȳ��mB����-�8>�W���?� ��'w��H\��������i�������=Åu�4��(�ʠ�?�6�%�<=�	j��0z�A I:m8�"�9C���+ת�ia�I���e�i ";�5*��t��ˌ��'��V"L���V�����'�=<Xv���>�aA]B��B�J��r��I4�\���V��%(��'H���_A��4.�y_��L��<橅#Mu�  ���W�{�gQQ?�;P�;�!y l8���88�8������[��dxH|'�[a�ּѹmg콷�~ >���yۮ�-奛�oW�b�j��tq��(]>(@����iӯqw�0�ܲ�O��*&#dRP22LpSO��_����$����#Z(��ُ���X�����Qp�����CC(� ꂾ��h}�c�Ys'������}�Fp|̍��*��jW]��x��h\dk1[�-�L �x��������_r�s���BV]%�>����s�̛6l}�-�`�t�����=?Z^�"���0α~�M}����	%��G&��Y��E��j��@o�9R��V��9�s�����J(�V�Cb�]h[�cG&����B��#��c��uѲ��FM%H�f%�*Ψ�=��T6O�As1���ʤ��qh��S�W�<Q�fڲ�f�d�����=�������Dj�␭,-�A	Oe�����o,Y�Cr���!��و�2�s��N?G���(�A`���~!Ԡ/>@�oS���j?���t;�:���=���&�l��Z�/1�P�>�7�P�Lp��~&�E����'�Yޣ����@�K ��`�9���"%������_R��c�/-#A����݂Z�ܶ���Kd;����
��!�d��d뮊{N;�3U΂V\Z*��YR����<� � ��!�v/y#R��O�J�I��g��qe�Tq�Ļ��&��7��6Ü0?�a�ZW.G̓�n��AQʤ��
Z���V�`=�:y�9��A��DD��CB8������Ѐ��XU��?)��#�
~+��Z��f���AP%j(sV���4�ǣv�5P��:8���w;03k�T���cte�m����9���J�����M���-f;��2Fp&�3\_��('N�@�����a�����e0	+/~���l�� �	����l��r�NR~D�(�4�ht<_I�f�6�j��"=t�:�����F�l^����-�xf]nQ/K.4-����� v�F�"��4Z�p�p��5�` s�F:�^д�,�}���x��'�<+�G-�7�Ư3���=�D�%����5�^s��{V�w��/Q�D��h����_�a,�'s�&�/�����R�Np%a��0�/hO)�HAy�V�txQ��d[2C�{P��L��&�ᐎR��q�L������]C�8��]Dx�) �%�W��*S	l�Q$���=�%�e�����x���j�{�[�Y4�O�R�Tz�Z+_���dZлii���努BY�#	�	HJ�6#m�Ç�4[^xM�� ��J��9޺�)�43T��7�6�W<9�n��5����Ӹn�?�:�8�Ny���n�Ćk���A��~Ĺv��_/jƀ��/���%��\���r�eeR�#���a.���r�L�̦�W��^�͈{�����N5'T�l��T�Q�H�!�
{@�&�kh���ŋ�&d�\�Gć��x ��'����6��;��C�~�t��Q^��(��3I�B�P�w�.���[.�L�V�� t����?uW8�/5������l^�'-8�����9��2�4nO�.�Kpg��3^�@�T��x�X�<o�
�"��Fh��+�9��,�ry&���"�ƴ�<V��r�mk��+t�Ӵ���0N�A��;��0������|BN>��u��^��v�(��Zf��F������U1���q׺%6e'C��@Z�H��O�h<���)U�_[ގP���Q��L9�Y�9N�^���5���*[|���M�-�@���x�F���jJ.Ӿ�m�XB����o�./dcl1��?�y�9�u���?+ՠ��F���}b(��Pl�K��Wm0����/�t�-����U��R�Pn