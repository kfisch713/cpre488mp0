XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��P���⃣�	08��G���/C�D&��A,Ah�޵)t2aA�S�&Y�L��BM�0�8�0�����&B�~�r6�?�%��jO�L�e�����U�ˎ���E�CK&��ϟ(a�*�'J� �TȞ�N��+0�l6����q����p!F��`%U�[Oދc��l���bb.��7�yn"�����R�}��riݕ$`d�1y��1�����Z9�k�Ԯ6����/˖�c"��
��
�Lw�"����m��Y'�@F�����%����~� 쌏�#}	�X|�A*��'�rw���� /v�^H���iSRs|���+R	���̃�E�H̛�7��0vz��b��H�����^+����o6�}.���S�)߀�~��)Qm<�4!h�A�ǜ�?�,����hJ�e�n���*� `T�flA�f�r��B�?6�6Y�[U��~�+���)Ԓ'NOk&�{�=�r{~�?�򘎟\B��J���i�|�/��}�y�p|���C� -Ph���6eۮ�W�l�����A���uLj����*]9V��yd�qx+&���'}��x̍��#&�3����y���O�VO�����a{�_�L��{�-�����	����4�'ӏQ��S̜�fyK��.�!�	k�W2��F,��<I�<�e�/����a�6�s�l��D0g�{�,�M��W8��R��r�u� ��A ���"�2��4�B�U�<)�Zߧ؅IqF���(�-�o���XlxVHYEB    1853     810�˘��A��[nS�֫�F%���[S�ܟf�a���Һ9NO�3�B�C���D"�Z���ԍ�h�����3�dg̿g��,}�Ʒ����o{,ei�� ���0�7g	T�����*Bs��'��{��g�	ɔRZ˕��.FҲz"��6�#�kX���T�vvvN]��K��.);��y7���(X=� �I����+V�m���9����Z����W��DI-���r#���ҩPX���ǋ��+*�s��r(�z��U�:���%?]ݡ͂$�N��ZV�DcD)+�Wk���j�&��Y=��	Q�/���2��Hyh��8I_{%W_��k_H&�����~B��HD���6�O��D��I�K�:Z�}D2~����k<��� 	(��\��&m,Ϲ���-�a�3߹i2��ӕ����V��[)��P��mBn'p~��p�|$��n�oW�*D��/_�^A�{8�4;�Y۝z�����">1�NEG.qRPS�׫�רe0o�=6����Y���.�Zd�·�ݮ��Q8E=v�_�w���!S�X��K������)��y��2�U.wP��Fj�����%nl����<�DA���Kzcr�^�� *F`+*Ķ���9@�� �{�^3����8I"�FPI�d�ZM�c����>LR�w��iZ�=ceO��������-�;��JB�.��-���6��Tm��~R�}Y�>]pv�#�
.�%��n$N�&�4qV��B/v��@=W�� ��@����Pg+�A`�-��A^���lk~�@��O�
[kIQ~�B���?F�bǽ��
WS-�[�}��'SI�FD8| ��h>i�e�� @f�k�.��z��YM�om)Q�eZ���Z�3W[-$s�����0�(,�0���?H2z��E��z�j��OQ�_Q)�6Qs�l2c^���]��G7 1���46���dJ���+	�@=0����~�X�E��y�en*��!1�]��1|�'�{��P����n���E����]��?�V}��ue"������WH#7�T���4�m�2~`�}��q�ƛBv�d��&7�o>��l6Px�*��ʗ料�G߫�vb�S�[�x%�r�ft<7+��U̦�`Z��OF��wab�a��|sи��5-��!��ՙ����Ƽ(�� ���7}�\�5�<���<�%t����}ϧ�SƄG����'?B���0I�߈O��A�ʱ�63�aS�fO�wv�2/D)Y�tȭ��x�/��f�/�~�2�i�~��3����I<:�+2d9d�ɬ��f��m�ġ���VCb��e���/��kn��S�>u�Xw�_�X�@�?xE���Z�U�́L�
�S��<�k���~�k��z$e��<�:�����)�V��Va������)��{���(�e��@�C]W�}U"4�#�3�x��YDrOU*ɧ��&��I��!ap�3�;�6�Ԥ/.�{kM��z����%��E��v�}E���A����]@�%���Ig� �F�m�5��َ�0�`���(�Y�p���cAP.��C� ��Wη?�v��zs;���|�$ȱ��=\���D']$�"���"�� ���I����Yfk���x�p�U���O�R��K�]�(�@���t1�U��n��@6�<i{*�p]�ATv^"X��vy��i���)��t�����CH"!���B+�H�Ve>{�:���S�3��Y��ȏ�Bq��H?�g$�uA�O<�<����^����.$gD��d�>K4���K�c�ěpQu߉(.6��|��&+W4�9�]d�}���@$�nQ�Lf��L��/�CTu\K�DMk��j��2κv*+�������)G��\v�#��:u��7�ơ$�F���<n�G�c[@��^�o���Ϩ>җ`W6f�
�gI��/���[ȏm�����'}�!����H��a
L7�P=���`�N��<{���x
�f�"+�P([��0jX,p4�l�J�>�=�o#'�ܥ9��