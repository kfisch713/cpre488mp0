XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���m��K�|#�$�,�vIh@���?�BvEL�"��o�8��Ĺp�8OoT�R���x�o�_	���Lu$2�r\�s�4�%��r�B$Ӛ�KD
>���z
p�3s�D>�p��J
��E�JJ���D��r��'GF �x�"Rҩ�s�:9�]�����5�P
��N����ԁ�Լ�]��U�z�lR�����-S��_t��v�W�Vˬ�	f���MN�<��˳b�E���k)+I(�B㷪�j�ń����S�~椚�����yz'p�[�C+�J�=��ր���9DC�5W���qc\Jݍ�݁�Fs1�JSd����h���f����z��V{Wg�&�5��`�[aK2�(Tà$}�7��i���J���ّ���+�m{*��3������[��u���L����������E��h^~�sLCz�S�߃�L����f�Z3�/��B�J��I��o��f���e^^�q>l�����]	X�ʀmi�����L�`�NMBLú�R`��#n9���[��f�&�̎�+��B�c�K}��o?�P�� �f��>�0 �\���j�r�d���y��߽��=�ܑ44���c��n��4��􍡟iY��%���؍����#�����D�G��O����.�vN��/�lڷ|�G/�/&_C��,��A١�;�Fu*`b6���@���,��km�Ѧ8#4�Z��H���Ro|����g��'�� �;t
qNJ�T1� y����>��q�c�Œ�XlxVHYEB    6014    1840(��~�`���#��!wG�!%�֥s�M�C%<ԯ�e���ŐQӲ������F�W�K��[�ʧ�1�koT@�'`��$⿽~��%�I�e,�8��}X�tW=q��z��7�N<�H���Dދ-��8��M��������YR�͚�#����q�gڃBt/h>{��M�|~	�=9�[C���9�5� ۜϭ��U�($mM��cf '�ew��`��#_�h�;3�b`�)��b��l�r���c�p�]�����o�}"���0���#_/j�s�tX���f�ϔ9��]R�Q��r��OF����g;��+�sg���c�eV�z�� ���4�rچ7٣4U����e�b	��V�#�n����^H�, �ի�>�61�U�f�kI�&����4i�}�h�J���k�M�~,��J�/�ڏ�@�Laɕ84{x(�g��%$�[�2wK%����j�H���y�������0f>�^O��g� ��?c��Hy��{V<�p՛ݐgJ�ݢ����"+��N�8�Ӊ�����{�wā�)��n��5��Q�q�6=���c�������"�+�]X�H�����d���dX�2�+��3��ƝQX4DWne��t��nY"al}���z�v&��de��쎲��U0~n	]:�OAL�� �����Q>�BGN��(BH?��w��n������)^ƦfhQ#Y�Z1�j̑��{~~�#γ����u�첥���dĭ�/:��)�x�,`�}��VN�%qm�w�m��^��Q�s��3q�o0�:'�/��1
�京%?�E��U�Fsj*��?�P���(�{��XMI	扊f��jC�F)��Me���+F��M�����SX��I�l.���lE"�A.���q�^P�	�TxС6_C������Gһ���<��^����Lu��	�#$.��z�zC���)HHX(��*5�b=��M_�T�߹B�<������s��["^����i���~I���,Y�cH+���'�	Bq��؊E�̎��7}��W�+�<�y����U�>���K�����ʩEo��.M��W���qeD=�VWo��8�-yl*�� ��4���z�:�<W�$���5�EmW�,��2J��RX�B'YD]��a�j7��� Y�䗠���&��^��bCy���n`�L��E�Xٯ/@c�b7.Z���/���AZ�H~6_P��"�M�+��:U&�w��&j &�`V������4�b��{9pyS��jM��n�V�����&,��� %l���h��$L�h��	;��<{_��n�[���Հ��.�o�د����|�ڨg4#��[�ep2p��}֨���guھ�]D}֎¼[�/����{E/^���D�6g����Yr{��B	=�2��4��K���ς��t=���X^��kX^ߏ���0��_g9Z$F�0s�\O��K��b	0_�'��@���uq?���4Y�A£IO�·�	��q� u�g�_���*���!]�o�˭]�{p�l��;�__SV��b��8���y�.�7�ۈ2?�A���a)���j�w��#�;=���R>٧��� ��z�5��%��#,+2���N|) �v AW��WvTR�9�������%f]���9���H��Lu�K⏞�ۙOy������BGU�8��@������n�s���)�PN��a�[���_d�l�~��Ll�#���(a� P�0pْ�����ۺ���TsN��3r̿,"Q�n����A(�J��ǋ9���IK�֨��|ʋ��ݵ��)��j�X9�̍	�|�� � �KR�c�,液��c-\�{�3�)�Ui m��n�Z#{D'��T�l�����loO��y��7a%��:^I�\5�ث驺zgDfM@h�ؽf�f�	O�G�����*C��I��sc;h��>6x�4gf~���5��'.��c�F�1���ͣwj�[��w�ۙk�*/���E�
���Ze����*m7��b�~[�_O�	˦����Ȉ�/��D�#��4��о.]����D���۵u�lsT�	=����+��A������&ؤ��_� P.#7Ѵ�qn�t���e�~;����Rɇդ=j����w����:y����P_5/���;T������
��v������ڌ_��0���9"d�N��#yG�(��M,��_��9�+��Z���-��X��?yU��+?Siq=��s�	Ri�{��y Ӿ��5o��M�xEv�����*���y�/����{ ��K.%��'i���'ȖƳ�rL4V�q�k���o ���5�=�P���U����.5��g�,V��kyܜ��5�q��75�����t�ͭ���G=�E=H?�D:�����ϻ�����z)N���X"̠����̝�� v#�{�֢��E�t��T�����������7��ZfXO���6�g�Xf��x���J���W�4�ik���>B�I%���_{h�&����A�PO�X
;wOx(~�6x-F~�,9+/�ُ�w�Ў��s�ϩ����ǣ9y�S�y	!j����7^�� �=�\U�8"zc��S�j/�#0��#��6a�Q�C�l��e�E���`�S)e׆�1Wե�����d���Tat�/�+�<z���Z�K̢Ï�� 0����y(��T��.R�}_RL���'��>d'�er�m�B��b
� M����S-�����oGX2O2^�,��Y.��<���ng#?�Wf����uv(s�l�B�b�{���vD#�@���Hz�^���]1\�q'�zJ�(��b��ظ�~����?h��D�򋨱e&�ۍ��P��t��+�5Y~���I��F���\�C��6���6@�oJ5ԇV���"�P
~p?�[�� w}������/G5͸��H�F�f��z5S����k�}Y�Jroy�ݹ�����D���<v׍��.mͨ������X�&��A�U�� �W���Ё�f��ͽ%L�?�2I���>͉��J�1�J�����Ճ��
�%�f���.���u9|�gϾ @4��1[ c/��q��*g�5��}8�G��N߅9�N��/!�0���5i�X�\�Ǵ�'��M�ɸ��Y�q7�$� d���� �
[乲m����m��l�����x�4�8��.��ad9X{��t�^�K��a�'�7�:�AߘUH�kqEMF���#gL�V�ɮQ����,ޝ!\Y9��p���f�P`�����݌��e�XE�j��mg��>�cϽ��H��7��H���� R��?r`$Y�z!�T�yX�e_zs�֙B2G�I�j�|ʧS���e�W��;}�Lju�@p�-"�⻃v�]�"Rn�>��2	21vi�UԈ�#����ǣ*М^�1p�w0�l9&�d��!����d���N.rH�DU>u��	%ݦnd	�������Y��h��r��*j;��ϊw�B���G��KQ��.حT��@�[�m��#v��+&Z�jc��H�y�@(�*VeW�S>G��1Q#6\p�SjI�rl�~Vn���nx
���M�k� �*��0u�$\"R�����KV�	��3NtkP�~�s���v�i���;�ᱛ����h$ol�n�C!��"۷ԙ��_*`�ϑ!�'n�)*���$�����W�?2˨�֕A��
�3�^���-�My�!�j+��n_��;�	���pSs7���Q�ː�j�W,yr�G"J�SDq9)�W�/%^uI��%	�Ƚxޅ��mB���/wy�V(�t�F�������$�N2��M0�u��cQ�Z�mwx�L���S����S��`m<��U�M�A�����P?��&�'���Ņ[�q�1L���d��Y>�;ު�\p��,&�9���td6�m���Y��\�ITz��AC�Qz��CM�<�:�4��R���9���{�04׵�)�u �k_��c�H3gb/d*�
�x���[�Zr>>�.P*,���x�D2T|X��<�q�6��7�ғՎ���j>NQ�Ih��7D�`�cIM��Eᡅ2�pK�+O�1Z��YG�FQ����?��&��F�(tc�R/ʸ�oP����'�S�< glo��x+�
���������G���i�p��,R�֠ᯤi�3F|s��	\^��;�c��)H6�c~(���.�/��R~8a��ꣶ����+8I�T���O8��w�{D�e����s�?��V��U�}0a��@��� �<��HxWP�
"T�53g���`�b��ݲ[]	OHn�W��F�`3��2z} BtR�����\��::=k��]L7��*�� <�@��){���֦��r�a&'p1���,��*d�5gG7��P�}�*�[o[0�n2�V�L��M(����Er+�Z��5j�ȸG��T�7��뚆⏋'W���C��6�M����n=}5��>2C2�}	z���$�C�Ե#SY��U��`5�}8_O�
�S���Y����	]�厱Иi/��Of5^��@�H�#�R�N�Y�ہt��jٶ_�|D�<ĐT��� �����w�z��p��~I��II�Ҽ�l������jO���ISt��IdÍ)'��M}C8A�j���R��DTQ��lV�0 k( 4�hf�-�!o���T0�<���¥yqx;ݶ,�� {#}2�����f��i���X$|%x����*J�*��[���c�����R3o/�� �cC�}�9$���qL���a!e�P�H�Frڏ�|6H\�!�H�MO��jw�.FYmy���r�����ً���TƮcPh\t�>R�/�v^��-��$s�Zp���,�;@ڂ�� �,'�/����2m7̍�1�y��z����1&D� �B���V�8OD�81�"��O��FĿS ti�1�2��q��>?��/�ce��cs|U"��?��u�{H���J����f*د�琶�g��չ��f~��`�w������0�Q���Ù�(7!�����@<�l�@y��R{����T}�e�j]v'�N���x�D�	#P��O\���C�n(L�U?~T!}4h[�х��Ȏ�}	=��+���Mj|	��%/�*�$ S�O��礠�߭�r-��	
�����5	��Ӿ���Eb������:��G}��\'�Q�l��$Ք
��j~�|�]��%�7$(;Ǝ�:�x�[֩e$�W)u���T��'3O����gn��_E�?�hһs��5A�u<����ݪ���&��l�����Ƿ�Tٵu����&7Vz�����̵<��'�_���*��X0R�Nك��C~P�������*�,���va�cc���ui/��&K)O�!���q����:���_^)���V\���^URhJ,i�8ќ�G��&�($k�-W����\�E֨$��l�������Lh!��&��9f!墫���dx���'��T�K�-���Fַa"t�b�1]��dO��]8��i�� �{�g�;�Y�l(��iR�m�R<H5��S�=��p�X�?GCQ&��Ŀ~�koC�M��A2wmw�+�X���Ç���t��Ն=�1�)&�h	c)/b5��@5HN��/-a�J��2����}%Ҳ����B !x��B�T����4��Q��յ�%���zX�$AwhQ+��v���g_7P���u8��,U���[�568r
<+�~��G�Q;���bqQ�S���@�K���j<I'Mca�����@&��]z*�B���)��+�~g�2�M��Θ�2�q��g�餿U9�#����R��{t���I�|5�����^Ě1j�I�')�l!Nd r$�tJ�0��0G�Œ�c�F��h�"�|���" Y���BBY_|��؂���e�ʕ�>�>�ƃc�\�w�B�2U)���a<� ��-��I������l��XūC�/h���d��P��Y�n3Ӕ�'D2���ǲKF���mD�4�B�Q�3s�d������1�7^����
ˈF@1�I�/��V�^~��ߊ�=�����,H�