XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"��
.��+����f+mG�~�<lҷ�t����&�-�Ż<�ۯ''5U�� U�Ro�Y`>���RC����L�0��})�-
&��� H&�:�R�dl�
�d�7�1��7"��N������6��?�<��M$|F!�'�#>�	F/��ŭ�:7N�Կ���7�C�?��g�:8��x~���:ޮ����/x�r��u!�-�]��j����.�°�t*��|iu��/���E�u3�f�Q����
�2@�4�r���J&'����#&T���A��C�����+��N�P����z��� %n�#t�=�b֍aR�]Z�x�]�wwW	���>o-�K{j�9�SP΢l<]��;�͙E��̐�ckkf�Y�Fٝ�� �\U;(-E�P�"p��W�Ĉ����kw��w)r���r|��pDZ�Q)s�^��YE�5
��y���'����oIh8�Hz�N�]�{4�����`��ր���r�"$�����P%HQU@����<>.�`2��p�ƞH�	-�>�t��.�v�5�d���\���BO�t��h��t���Z(�>q{O��Z3�x���C<W��NJ����~9�dӴ�w!X�Ey���B�+lY�g�nip�����~�,V�pW���Ǝ����3�V�|�嫉�Nܬld���G	�����i�P�C=D#XB"`�^�`�<���:_)���O�����5���_�0g]q~��)�{�s�>\;��П�&��XlxVHYEB    dd8f    2160�;�CJ ChdRt�g8��9�����S��tj'n��Lѹsy��������DǱ����pR�=tL)k���B�}k������!;RT��a�P��zP��{����`	U"4���$ J�n��]R���w�pK<\~�/�8rV��L9tBީ�d@0�*����s��w�ʃ��F��e7�D�B������K�V��BvW~�r�Fh�1kN�k�t�76����R���clj=�~GV���9X}q�Đ5V"<�M��u��$�V�?����j%qϑ14Q�s���r� k@9kՖ�2R<�3�tN9����؂�1t�e	��*�4�8{�6�Q�g��fN��N{d�6�����'Vf����k��j�Sѳ�下��N��M�n�G#�cW��k���r2�0�Oq�L��	�����5�'[$�����9���q�ԏq�[�jU)l%�U�P5.�)/Ջ=V�?ۻ��:[��T�0�Y�F�I�iD�@�����/?
߮L~5��/�l�ot�L3�:�K�lU.`�\e�Gm|�]���2��K�����퍞����7�A�.���g�&hj��"�.�?o�ݟС�R1��,*}�?���uh`W
%�f�X @��=����N�n!?]��~��P8�&�F�uu��N1��g�e(C��SV��'値J��� gq�ә�{�C��r�]mdJ��`x���؆O�G:�-ɞ�j�٤���h��ߋ''�����[���H��<�EC��W���8�;��¡l�����l_c�B���G�y���y��Q/�j�5R�d����[�N`s�W��]tkW�M��<�J���!BB�� ^��'2�0�W���2z�c��^�|�Y��;e�"«X<��Y`����Ɔ-,S(#� �ŭ����+b�����զ�M���[ҋ�_;P�"ЊMD�5�YUis?h�{d35�	|䌪"��i�(�a��A���`��چ9�Q0��W{�_Yy]�3��q�z����yĐCn����y~PR��A���|V'^����i��p���m�$�!	uerq��_Q!c_#�a~=�+n�7?��S��cT�ny``dâ_�J�ۺ>JN������Z1~M�I@17c6Ć�3�ބ`�J��Uz|��V0�4PK�� [���U�c�.��r���tG{ܠu\	���P�ge\���;`ƥ�+l$�eQ�Ń���ǂ��vG효|���L�&�W�"�a�.U�=Ob�F ��k��̟k{�]��k��=�PXqI)rEsģ�6�A`)���$�� �5(��ø ?�&3[�]\�Y�N���=yz{X~�d�F�	�j�b�Oƻ�\PۉBq"�
"�9�s$8!4�g���(�!���ݢ���5��1�W��]C�]@X�\����F��J"������0��R{��t n��Et\��$��)��@e)��2a5���I	jQNz-}g|X[?�y���z�Y{�G>-+������-[t�V��0�4��$A\��M��x*�Y�ޓ\�_�O[f�:[�y�a-�����bg�c�}��pܸ#؈�\߫����n_1�D�ֳ�����X�P�?�1�����ہc�zi� �t��k����(�X�����y�-{a!�N�O?����=a���M#�9���E���Xo����g���A�&��k�dXH�U�f́��TY��J�p�\�\�&��_uu���C�4���������)����P�%vw���/�y���tw
�jf��C9'kGk-�Y�Rt�Dp�Z7JYlm;�߅��<6i�5bwW�[�m���8�Nd�]��h�-'j{���s;�W�9��2�0x��4yD8+U裛U�C��ԃ��	�$��P�vn�-_�r�SF��]�B����nC�Z����00-�ئ$��/D���=�~���kr���H��v�i�:��(��A�JL�>騸��OGD�*��tE�_�er��Mm�U���|e-��o�dăF�jfr��4��֭����~�7]����ʛ9j杔���dϋd\�,LA"�G��ʢ�R����~v��v��Ѕ̣�)�L�m�h"��u ��,��
���p��
�Ϝ�]|�uC�T��94\|�'��?R�p{��K�1�H���M$T���W\�H(���-��@�c�Nv��re3��0Hfd(�tF����F�U"�[�+a�.?��3'�k������Z�x^*�����p��w�R����rD�?���X�[��QV
��Nt��!s=L9���Sg��~������O@���L��V s��n����'���F���=���z{~	bB��%y�n� ٤U��q�Y0c�Y��y�`4��V����ů� &^�%�ܼ���G^�("N�t�z8ղ�w޺������fǊ�mR��M�FX��Q�LĬ�G�lY㫪I��,q$�b��Ћf��j��2I�.'h��?Lw��9F���@�:m�P&���@fh���k�6笰��{������S��nV�Cb����zQ/���P���Pt���tM��XB��e��&�Ҕ�ֆ*B�R��'�m�@��M����h�]F5K���1H�0R�f.Ϊ8�ў)P�dl�6g�m�4��ټ��'����1w t VI|��2	�%FRRѡ?b���n�L�s�HkU�s��I�.y�:�Ӟ�u���đup�|�:������ ����K��ߐ��l�3�+�pKC5�s��Ĵ��� �nI���B�����{~���1*O{��v��y{����L�*��[Oh��o��F�Xqz@th�z��JFCq]q['�lpK��q�� �o9��-	:n$����͢�z�2����������׺π�Z՛�����F9tS?l���%�-ќ�Ĵ!����@ks]'Ο�_ �l�#<����������h,ܯՙ1
[��L�!7���a�Q��ߗ�f�3Ej���c�Ɍ�F�[GgCUHM���<:�q��L��q��e��_q�kI��9�I�I����õʍ�o��ɸ��Kd�3��Ȑ�2������/2��|sz\�1(�3�a��@�8ٹ��W��vc�ܲ:��04���D3��D��繫ݏ��H̺\�tح,L�[3�:��� ���F�It[,�Ҡ�nø�0��2�][v.���u1 �0=}#����!/��q���잗q4�h�i虜�=K�����0��Svi��ʺ�Σ2r�L;m��q���/
��c�␻��^��к-���e�+#�^�+��Vy��f	�y5� KGo���r^&��~��������b̤:���g���-Y�A�s�=x]Z"��Sh�,�%F�o7�����PB����������v�����_�� *e�m�o6��Z{��{Q�iY*e(G��;���Pg"�z4�WWC������ʭ�u��W���Z�t1/�T[��x�<�P����(�G߱_��22X1���^3	T+Ş-w��ݻ�����WG;�uxjqa>i�����x�Q���t�Fr�X�؞�D<�5g���������L,��(��E����b�4W��G����.�������|�R�u���]�x1��*ޟ���K�`��k���j.z^�w�4@=~� )�Ɇc"�$h5���K�b��g8mв���RX�C�`�4�����-b<f�p�%0xn���Fn �-4��e]:U+�~��`���a���:��v�����"��2��N������>F�Zۉ��T�:_
���ʙonB��#�k��b��IIz��~�9#� �����ͤGW;ò�S`�?�������(ԫ��,���"ԙ	���0�:1�f%���9��SF�ߋA���?ѫ��΁��B-��VC7� HRu��Mj�Ⱦ����+.�ݧ���s�_�Q��v텘�N�$0vi��"��zL���В�%^��S�U|�^`y:�����	�5~c�G<���(�s
ð#=vX[���(@�[�0x�^5��7�
b X�&;���H����jv!k��0���vե��{v@��h�����qqnЅ����Up���Q���f�YȄ��A���>�}��_ 5��^"��cT��qsE�D�X����7�A���`O�#�s������7E5��V�c����f�� �t�[k�r2 � �#�peN�֭��,k�H������-G���'�)���w�WP�zUћ�8���P�ǚ@�l%���q8 �� ҈-�<�ڛ=��Xc�J�gf�=z��XE(�������˓��!T��VH�`g߆ͯ.���M:��^-J����`maa�<�x2�_�����PR!�;����<_&>I|�?V��G��'I�HB#�����^���rT����r?S�ʲ.�Y z,w���ܲ��w�
%ce�
�IN]m��8�}�h�CǴ�'v7��S���H�FH��ꈮ���ȝ 4R���h� ����o`�23�r�C,Lc��x��n bK�Y�ȟ�� ��:�b�}�+�$��8�b��h��V���m#�("�S��GW��+��H��d��i5�M��BES/A�����*@��������uqT�2�G�}���W�4�TтHd#�
�J7^�%�� ��Y�9]d�*u���>�ZN���<��D�f(hN��7������iLx&b[���tYZ�PJE�
��R6ߒ,1� �>*��>#�l?�k�D�L+��U�*ԝ\ϐB�"�k��BǓ��msZ���
Նxr�R�x�&q2���ߪ����R�k�ۄ�!q�aX�Q���l?�3��Хț����>Y���� ��H<꯾	�����ݣ��(NsMA)�y��E��tNBd�2�y֝�R3���&��{���/����7t��$I��G���滛���EpkD\D�S�I1�0�A5U)�u�,}'�՚����4V��sqI���&�DXZ}6����8��*��qUT.�E��x�V��D���%���^{)��G�9�@�mL!��~��o��lXL�w�0,1�Jc;l��gGF�E���+'��XO���_��ܧ�$W��p7c���)�lͻA@��,YxwVk�T�o�!j���h����=#���V���,A����i���?�c�,��
z²3̌c��S�P�4.Tv~���`��|r�h�������M�`�h�4��ـ!��|��
s�e�+�6:�S1�f� #�j��zDN��1]Hm����H�C���|���x�&ߗ�����F6l(�&J�p�~��*�eo�j:����O��@X�bQ7��w����^�O�M]�g@N���U��X�T�)iEK�/�*��s^n���ab�(&\����z�%*ē���B9ḍ�M��U�rh�yf��D����У-�1G�j=�D�Ճ��\֭P�PO�����aU՟B��@W��,%m�/�9d����U�'��&�_U�?>�3��^���-p���<�F���#I��}�!��h��D��X�R%��i�_ߡ8Y��`�MF��t2<���.��T~�d��ξ��J����j��]p��mT�5��mjn'��yǡA< XΕ���E��V6���E�� �� x�X�2��%3��Pr
S ��$�w�p_z��E�v�$��9�X�'�� ����	�� �� � c��_��^�t���B���=H�fŎ��mp��<-j��@S�Ez<&^��+oJ!^�7^�F߈���v���l>����Ԋ%8-g��d�5	h���:ȝ��e>|3Ř�q��hD�Q|���u�J֤(x�
K+<�M���4fˌä�K6���T��VS�l��]	����p�Wm+��iMi>�T�*uX�Io�tOM�F��`��!"/[X�O���J�����z)�s��e��������84�3==�}����6�!�<J��_�N��9�H��á�2��(ܫ�{��m��MJ�X�5M�����8����9(U%�NkMG��ṫ%]�se���@�`a��&�П��[�Z�I�I�n2�w���f�
�UE��=X���r��x���5�C]�r�Ȅ�L�f1��/ƴ
&���ݺ1B]V�Y��a�9WX��Pt�e��&]�`h�Z��մ<a�23	�����ߪ�[ʀ�8C��N�b����=y����A�����جq�&��!�i�.�'U`����E������&�X�_�B��� �P��7z0i;�wʮ���bK-�YQ.��U�v}U*��,�k�і]�|k���tl��m�T?H=\c���1��k�i�l�S� ��];ԑU��gHû?�m9�Ep�GT>���h�FPF��`��U�w��  ��d7H\U{H��&�Og�y��sC)⢆��t�?z�����R��T毪����>�60�Ҁ�v
��l�sW����~N�j�c���d 9P�v1	Pv��F���>���@��x�ϼ�u
wL��z��T��L~��-���$�-�>.�JoNR� �7�f����"�sc�A\�î㑄 ��<ufF��sq����q@ ���B�Y\�uZ���޻���!t��U���E#�gգ�*Տn��}���*� �_@�&-��-2 0v�Y��K����}�T���OUh(:V�
�vW�8�ni�2�Q�c7ּI^��fv��qy�\]����J���[$V�U�p��h��S���?�/�XR��+�{N�S��YI�ؼ���p/��-��D��ȑT)Ե�ػ���y��b�Q�q�8ԞԌ>!} 5�"\	�E�R�t�;�u��6�L"����A�:j��y�#ƣ���q�[��a�Du���?/>�Վ�}-�P�D�1�	��Q_w-�.���N��q�qE�yb���@�.�}���5 fI�O�E"���υy��f�����X6��2��꽿7�}�=��aQs�,'�ZN��لR'��bZ/�#V�6˻�O�1�NSv'�n�n~Z��fW���lf`ҧ���_�����Y�^��h{:��
L |�K���5h���Q�Ӓ�,��q�|o������:3)��R\������7�d�.��m-lی:�j�Q]f�-�u��6f���H|�V���F�O'p�j!KP'��_$�T���s�)�q�ly��T��>H�=qQI�1:��=.��oo�=pV�b�������|*�l��.Y����D1��pޣ�rѰ��N/��
E��7[���/"G�z{���� �+��1M�5���J����
s�7;-*~n���#J��([�����\��M�rdBnr��� >��4�+��R�.�?+�kC��� �d�%1?��SI8P���zE��q�������s���-M��a�	G��)Ru[u!�4�F�O Q�㮠mMXv\�R���Z��(�? �Ft��JN)4��ת�{q�β2`�Up}��S�42��){�k�o�w~|D��B�'�?�A����|Zx�t�n�#�S�*��o~ZoĬ��3Ṟ$�S��c۾�����浧����1�i_�-�f>O�'��J�5N1:"�"/R&��qrDs���c����+~ �NPP�ݳ���)(��M���{�î{KV(=|�2����^O�b2c�Q�5v5S�=E����uA3�B�GEg�ĵ������������1�@�v͵#��j]�-�������N3n�K]5E8J��j��Vx��f��{"I�R��Q�o�ɥ��׌���� B!��
�դ��� ��p����t������1�$j��k������/���>����؊V�b�u�a1?i����	;$�X[��E����P�I�6�g����ǂ�u����i���6�b���B!H��n$����u%�k�/���\�Z�F>��O��!ZRt?hGU4���3Ef)�d��ㄇt�0���jS8�Zi]�B�L�Z<�=�া��i�Z����5���R���,/��];OV`���EΘ�A!dN@rq���Y�ɵNiы�s(�::�a(���O��6g��/}	���n���J{xh���E��`�� �7ѴBp{��熸)�����PP"z�v��p��JA��a��7)��w'Z��ا³�rZz�R����v�O̺��ў@� �?�`k�@ޡ�����&�9u��_��!�;x�ݔ�a�ם�;���-�rD��Ү�ݞ�4I~Ϸ�8��*�;���SL����7�Zq�V)��D�El�rJ������ڢ�˶^	��89���țOw�v^��<����&�"�S���&����'���u�����;��Rdwxa���K��Ҥgu��Y,�[T���*������( swq�7��