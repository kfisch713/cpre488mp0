XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������e�c}2[x�i����y#%��$�z�a�%|^�B,/�*�<��<�i��h����;1��z���'�W��θ^��+"dml�{.�Ӏ�h�d,{E��Vq-��#$���+�6x�60'���"���A;��5[���,x%�qu-R%��^�v]�""	O��ff ���,�;Q��E�Д���'V�pˀ.�Y�e{��#/��^�E�0}9��
7��t�-1��m�Z\S�_�:��0B�}2�r0�.>�_BNX�c�x,b���S��j׾�7�Aq� �r���fj؅���r[�⏰��Ɋ�c����	m�q��>��޽��cL���߽^j$��9��|�2��1�)�A�-��B����`2�Br��/���_@!�G�
PD��R���g�P��pTKK��}���_��?s'K$���dt5a����#����N}��ޣ���֑P s�i�>EN�$��wV:�ͽ!ޑ�T
����;��6tŚ��MyaY���1���RC�϶�n�	�����DM���Rv���c���J���u�Ը�!L�z9�w˹��h�1p�W��S�Z^*� �qK�yر�	7�]x	�AY��c���1V�& 9ջ�����qKd{x��T��e�����_���8y�_��	��ړJ�������/�VR�Ln����<4���y*W���Z�It�&�s�{��;>C���wAD�g�6V���":��ID������c9�5K�Fy���XlxVHYEB    fa00    2040�"�_�T���F�v�L��O3t��?��%p����=��D��� 0Qk�qy�&���K�TN�^������t��Z���<����~�{���Y}'F��z�G���O%��P���p�H��Ͼe;�e����n��Tp�d�9�E��O��C�g6��<��}H���d&�uV4���|A:r$S� g��P�W큖(s�2)4��7��~:���A^`Ei3�S�it���3�&�� �^�r�ƣsc��0ݹ�R��vll����|�ȳ���*��&��<�U;$?;qF�|�^3��`��dmXG��l>�!yM��y�ws��x��\�S�*�.,�*<�C���&�&�\�yG0�n:�����ڙ��E�ڹ��љڿΌ�n�W�,�7]<Z?bv�O2O|C4����մk_:�nxj1?���ΰ��)�.�6�+�pu֩E{H��=+�Y���^v�pjܠI+a뚊��"  �f&�l���f��\'���y�q_����F�Cg܎�0)�»�3F�}���4�kr�٢�Pr���X���ô���	n�y���r��@��f�U���W3`O~%:�l�([���h��zw�b���\�����t����5���w޿G!�'%IM�hnG��9xw�(ôZ1O){P�{��
�"����jM�F��W�M�e��Q~�:a�*3*��jq\��@���z[޾��q,��$�8����1��p,n��|�8��yt���cf����!���N���,�״,S����k�UӲa赨}��k�ûVe����cJ� +�۟Ǥ�A�P�L������"M����0����؜�:�8^�kѭ+nX�o(�tR<�le��v��Јsۗ�����
.4�#iKۧ��/x�������S��h�G悹8C�y��t�� ����̜��g_]e��{h����yuFS��8Y�̺�:=o�}�L*��-M�F��-��E�/��Pp9�6MH{��w0���b�������%���y2�+��&����u'l�l�pm�Ӏ܃o��)�_޴!�����W�f��xD:����^�����R��yl�D*��9���
za���_�tbY�ept@�=�M�h���ֶ'.��+TvKە��.��*u�		�x����3ݕ4R:��(3�~t��+��ܷ�j��;t�5��ҭp���||�ҭ���NS|��u�|b��p6�wvڽj77���vX����U���o���D���J�Yt���-*�e��h�8�AC���yJ+���%�T ���z�U��ZZ���A�HgE��|�M]�~~T��e�K������o��Kb亇H[����w��I1�?P�5�hOvP��_H�c����f8�p�|k�J��L����X���H������X�De+.�of���S ��8A���!V�V��"T�r�kR�X�S��հ�ո����t��Bص_�(����[�~��qق��cҬ�F#I%�I���e�/}����b���૰��_�2��i)����E����gF(-fU��#��D�(��^�Fj�Q�ěN�uyns����V4C��Щ�b6	G��V�+����߽�H6 �i��^�OJ�y�χ��а�RT�@:���7�����?�+�e��xq4�g���N���W�)�ȅ�3_H�1���y��/�h��r=i�ջ;�"4����[�~�tBt�#����$��d��|�Ph�Jh ZJ?A��WZ��e\�\���8X(��|�6K�@�	�rK�e�&��2�����-�\�Gh��Ү�:d�-�v�N�T�>�b$�tM����:�I��p��v�<�(���Ś���1Z�;E�B�(���. ��N�&^�[N+4
�ቂp�k��ಆf�J���_�,��^S�4����r!����\�Otl�	P�3S6G��sp������\��8	6�I�99k��-l�� ,DN>PV�>��mx3��!6S^qL s�я�;h�̟�0��Bg��j�Q��"��������q��V�a���t	�5�M�܀Ց��5eS �fI�덡);^�b�.��9�&��?����;=D��wbQt��P @��.��X�����\��[��\7�-σy��/���s� X۳V��*�~�2n��� ��E��8ȽC���)P��_����7��i�@���4e7�զ�<�f[�x���-R�����6#
��u̅�,)�=������R�m��6�^�4��ԍ��/)�<��r���r�h��ܱ}	DH��4�!1p��v ��X�<"�����ϫ@8!���7�eP�?��{�&ϜY/�03��ּ���wp��f.\Q�:�;��h�����塐�ѯ��:]()�cHZC�eu��A	}��kdz=4C%�	t���Tk=7����
�}��a6'��P*�ʋ���"H�f���<���Y�����B�bHFj+�B~S�b����<��Ksv��[ʅ9�`����i��"p�}G`i���쑵`YAX�q�蚝��Mݰ�a��,���1D������Z�����#w�C��v2JY�"���M�8���pNWk�ZaH��Ȥ�<��袳��ǘs����(J�G�6L�UŦ%m�f��8����V�4g�"�zs�����<�͆����U�{�7�Ѯj8ock*a��4�����A���&�WS�1;����ǢP&W5C��4������+�/F�1�Q���/�w�w(��+v�(g�Q����)�h����Ĩ�ԑ������Ǎ.���By�o�C�O�KcP���/�jGS��*��£X�2�29q����'X%|����C�]!'C��L)������]J��1��M��V�՚�O��h�l���+�j\!I>咈���-@�:Cp���C����'Ϯ��#٨$'5п�v�.��[u<��oe�P�+�*An	�Q���lT�:F�����KIщ\�0�'��I��^�|(:�� >�x��XY'DRXv��릟k��Ԛ����܁r�q�4g���H7q�kAc���v[\1�����J�_(`����>�3�LE��,������F���<�N%�V���(R#}�"A?�O��4z��2�x?�p��u�t��ϻ*y����	�td�c��P-\G��%���.�=>��+8����/����"���t ��8�eظ�ϑ-p^�U���'/�ƪ�+*u�
��U���\�^�m>�@��b������`���E�-��{3��4URe|Z���ų��������������[r
�n$M�S6�S����� �dI������$�{1�ft��+x��2�E�YT��ۅ��NI��Z���|�������q��7,�K3�=��l��Y�^N`8�D�dg'����)1���fY���q�TI�nzyW��JquDJ�D��`,_��\��0��]��tm�&�3ֈ�r	C��5ѳ�Eʓ�ۺK��,@��������P�f���B�'\e�T���v	��6$���Vv�	�@�D���ol/^����p�X^�P���`x���O)9t�P�s%5�Nb�����%�0�t?$�y�a�^�x����^QXk��:a��Uڶ}��k6�-*��#/�K�T~�}�9,z0�r����M��a����uǤ���-@fG�R�(eI����0,al���#5� ��y�k2��=��ݘbp~�Q��_�i(�8���Cy�^f� �f� �A�O L	����.7h�Q����(x�:���nm�ù[P���=!�Ԫ`)!�9w�l�.�� 8�bx�,Ķ��ك}��\��33l��"��g[�Т�/hG�VV��:��b�W��Z�JC6�������&���#��Q�Zp�)�K�!~&[hCJU߬F������rr��� WG[�JdZ7��\���O��jdzC�Aac�3RY��4Cۑ�ܺȨW���!��-B�@���0��:Ya���1�YH��Dr%��l��6{O�&�C��*RtպM1|�i>	���i�*D�3z5��ŭA"�k��*��8�嫾��%r�%B6^oQ�"���?B���D����i��%��`|*��<I���g�Rߔ��8�Ȩb`<|`��t�Ϫ�`�,E������<�V�Tg�L.��+)�Wc�|cP�'��f�p���Γ��p�O
��ʝ�o��E�7���aݷ��,�<eIz�VQA=`���5�97����.l�6��+"���o��ej��N�k������B���7A-$	�y�a���|Y��`�h\@[0�Aj��Urbw�؄hA�����Aۦ�c8N&7B��>0d��8��I�{
M��ٹt<o������rA�S�4�+�k�S(��gILyx�Jg�!��e�u���m3�����'6h"B��m����ECug.&�X�_��!�K� �MA��x�c)����	T�<?j��w��O��]s�5	���6��� !'��$(����&|���g󁳾�~jK ,C l��}9갧�{�n��-�w֧���&�T�hE�K��������y���*�|��+k�J��f��K��--e�H��8���O�i_��ٖ8�7��qA�27P�!4v/o�:�GË��~{��F`�k��;�W���iC�Z�u�wr8�c!��u�p�d�&k��Yd��t��n���5��
���%8]i8��t`3��ZQ�7����Ò��&6����=6�����	'&R	S�_2���������z+*gTZ�����?��َ�~5~��&��q���w�W:\���
�cng���ŗ�&�1h��w̨�q-T&�8���W!�b�;�tp���h<A.�z�_�(��[\Lt���`����7���۹Җ�DQy�`�����ILc���# ����6�q�l�ku��v9�@MPŀ[ g�
4�����R�t_(7VSCeX�dF���1�t~�`r���?1�!
;�<���[G���<R���n�:ث�%�׷��h���z�� v�
��)��p�Xq�z��ɧ��j�hi����.4@�ނ��O�����E�o���^Н�a�D/��E0�($ .��L��G�������V�F����v�X�?x�I�@7Y�Z>�<rizs��r%�P��B赣�$A��8I��&���'vt�L���n��}e��;�pg�ီS��^I�?�mG�u'�"�I&�����^ș���r+�n6��É�B�w[�����e�	��@^��b)�p���(��g�s�W<u����	"�^��[�f䤈J����_��ơ�~��giX'PK�HKTbÚm˛�^J�j���m���DM�����^yI�N�����mR
�1"3q�k��7�b�x�/ 2���yU'Ȁŗ+����]cq9S�ţN���꙽p�!�Т��W臡n��#���N�5e\	�X�]�X$w�����5����o�L,Wo&E����mڀW5=u�d(���4C3����"Wm2�ٹ��p�^�N �i��Ⱥ"ց���}VD�#+Vt ���)��t�S�s�'ȁ��|��NW:Q<4MOfM��ȧ��XT�!���C�w���"Mx�S����gՓ(��!E�F���3X�Li��1��#n��9
>�/��#��)��mR�:� X�u�����4��jD��%1�LGH��H�`�ǩ!�zyA%��vl�d
I�0��X:�)�Y�a�K�֌�;�Y�T 6>T����k�k4���^�qZ�:�`���D]��i�c�x	�;
_�^�Kg�Q!���\�fؠ*Ygɖ냿f�qZچ�Ζ�$s�e���Kf�s����'+%����(�X7eQ[��n�Ԩ9S"\3���X�!�ҔB ;����qY��c��V���|���i^c���ޚ�������Ѐ�QR��<�JW�8P��J������0گ( �f���Z���.T^��s��{)��Z�H	_X-Ð��ouX�T������^���j�,A� }��9�"BY:"%��b�sa��a2&�=ǝjt<_�c7�9L�G��`f�^@�xn0��֘�6Q�z&����c:n��	�U�����T)�,u2�H�s}{���o��	9�5�JP��G���"�0s$�}.,K\\������`�r�x+���ϔփ�s��u)U�+s��>����J�&�2!��%�񊏺�,hĈ6Ƽ��h��5Y]-b�s��SJ��]�wb*��H��@���U�E��1�:�&�S���:M����a��	{��1��q����^P����j4?U�f�o#v�[�	����Շø����F�I�Q�4��E��<�e"��3�qW�"�ZJu|A�@�ڔ�Ո*�NT�'7�a-�`�����?�(#�(���uz�E|��=H�W"K��Q�C�uE���;�n�Jj@p��s����d����G�-qMǭ��ֲ�t*�U���X������ؐ(�Bbm)8| ���O�ڥ�̅}�=��C&a��S�Rޏ�)h/��m���4pz�vd��EB6K>���p1q�#d���(���4�,rYD$�e5�Q~��xv��Cl�W�;��1T�;[�;�M���ϲ�䁙\M����ձ ����C��6o�I��K�t�y�@Nq�8 C �{_�ʒ���~�|�qH
��"s�\W�Q/�ޠ�B-�>�-YjИO%dP�3��;o���c��8�Mt���v�#t^�/ w���]|h��/8��,p��
�>�Ъ�{V�q�e�?���P�����w�D�8� 
�64F&݀}��p2u�u����ZYŔtu`E������Z��=P��$>L���F�I��/iѴT�@�������'ʼ��1�t]�څ�ꦈ���#��6�/>��bĆ&rk}7�J�H��fP�#ٽ��*'�|YMVbT1�)R��rHQ�ef"헖�¼�i�W�C�C��K֧|�JM���d���l�
@��c�vo��N��ۏ83��nC0���)ng���I�n����,�(wHp�^����É�;Yk�k ��V��]���­�����K���ZP�c��y�@�D+بsN�+�jvA?KcB'g����s�x���h'�(�A�
���a�n*�ǘ҄�5V|���H���6���"<�ūF�1v�����ȍP��)@u)�u����e?�ӷcy�46?�
�d�������!L+Y&�z�鹲�z�g3��~&ԅ��3Տ��qg���)�m�l1y2#��[O{)���C����Q�0��?Nf��1XG��㗈���0�׎f�G ��Y�����C!��bW=W+5H�e�x�2D��z%	�ۓ&�g���4EW�4���>ܒ������_&�w�7���A��w̧�S
7���#B�������-��c~m�O�"en��,uǃοQ7xXJ�f�BHli��ǳ�y8�[��}��F�N��_"G�)���Ut�q/����<QE�|`�<�S�_�1�?%BL��U��#�L�ʉ]�'��o��k��T��j��y�#
��$�Z,RUØ8���Paɍ4G"pd[��ӓ�bwy�ʯ$�����>�����Yc�=��)���V�zZ�!���{?m�VB0���e+|��OR��d>��%��+q�i3�;�R�C?w=.h��%��O�	�N���m�㝤�i�.|{Z�U1�
qksj��V6��]�W���	���d:=k靳�v8M����0:�0��>��y.������ᬘ���ξ��1� ��!��?qd�z�,nRV�:�l�|߉���]�	�j�Fy6d�� 51Sd�7Z�Ʋ$� ȹQ�#p �\O���vφn0��:IN�����֔�8�PT�tłj��8i�&��ug��bDt��6�uG&���&�8�}�J��6��!U�C��]bo�/q}۹��0'�H�`;��#BL�c������7+���E���ޔ��%��./_2�jI�S�X�:�#i�Ex������р_����  �{X��f��O�ӥ�e���{��*FXlxVHYEB    4f62     b50�L��(�R:�>�F���HC>�(�n������pnJ��η�Gj��M �������%v��:v$n��Mz�Q��w�sl�w9y�E���A�
���9A��ii��!��y��P�b��g[5���6/���>���c��t��#����MI��6�,��2�8��q�8%O�q��1R,�.������W<u�]VA�F��r�ڐ���vg�~g���T�8#��h�l�{�C�>M:���X�1�׎��M8�|���M��Z��a��
�"����i��z�7%�l���l���V�E���[�^���f��d���Y�Z����;�;��}Ѧ���vu��Lx��s�0���Pw-�5�M�
/�G��(�+e�":QiG�v���P#a��t��f��Q�6�;^h�p��pYϽɔ��Z���{����p´q���Nf++$gi%�߸���A��T�R��6X�-�$@v\�bg4�
�o%&9fOG:Y��&�ⵑ�qI��@��;[�M�J��ew��Oe���s kgÕ>t�����N���!���]eу�G9<dW�����n��1D�R].���h)1[�{�s�̱�K����e5�4
���ޏ}7\��h��E�|��b�-�{'$����P;_���A��!���* �NH\��M��:�%׮�:V9�C��x�Ԅ�����:@�~=o�=�Zz�@d8�4��8��5��N�7���Ao�ΦA�;���'e��?)�~�l:�-A(�� �\;�F�UY��;ѣ��R�c1���U�������|L�g�]\�NEA�1��U����Xc���B�D�C������;�Qg��Ս�Y�W�P�A8�cF�\A:���.��=�"%e��ަ�jS}�-���:i���Fw�s�7F����Ti�u2���&�7�/�j�"(�Y_���7A��q�;�q\/�K������s��Y��pL�_����\��#N���Oΐ�5��{M'��T�up.��.�N�!^�	��K���f�9+��u=2�-�H,����_����KYk���J����!�ǰMLC�%�Fi�׶w�/Q�vZ�	u����e'/������=f{{�L���/�\� �N��<m83Fx
g��$b �ݾ_Ǳ�]����ƥ���wX��$���c|V�.�J��gH�KlUCt0�5��>��[=2�:��� ���2�4w�B�.�駈�+�9.f�p|��w�T�mVCu�r�H��"�(ׁy�_[��/��q�������&h�*tV2,���./��-�|�2��7Jx	g��9׆�[���W�y>�Y�9]��n�)c\<�c��~9���R��p܂��~���{�SV���&�g恃J1e&E�#M�DJF����!J��I��#��i�&/�~�8m��5��ϕ#�>/C&�ՒRt]�q��>m �Wa�o܍���ð.9+�K�p♈������I�}�_�ؠ�c	�Ϯ��D;�h�cXm�L�{7�Il4;�ó�8V�H��қ�~*w⧹��eAWX��n!I�:�+�`%�HUOo�M�3H�}:a�x����������o�R���k�+��<�����F֤�ֲ����ʮ����hV��&��j�&�+Y~I�!�4�ޟ�Q- %�(az�"ꀝ�]��/h�0��p=�(��R��#���ۣ�p�1�3]|T��I�[�"�X�L۩�χ��wf�g\E�F
��D��o��М`|��� ������EK��J���J�(�ܠꯟ̘-��{��n~C���w�@*T��G}q���hf5k�X.�[��Mx�3�*�P2A3}?e
z�~ᰵ���X�+��\�ڪz�W�O�ل"����r�'���Iu���'�Q����x�A1���w��>͈��T�_�0�b�ͫ�����Ed�r!��	6�˰��E褝��}��R�a���D�F�BkxOԾ�8�Gۋ�9_�֪�6Ϯ�ڋ.�e��Ź�a�����Y��o4����[��sR1�i?Aӻ�lj�W��1Dk��#��24$�.+ձ{c��e_���yl��C�2B�k�3:rm��i�%P>j�]&����9z�ēU��^[�`��#A�PD6c�B�OH��Pd�*�%�K�p��mˏ���o7Cx�����(�2t%�KO����Fқ�,��Vc�^r���Wx��S������A�0�~���J<�2e�S�}��/Ƨ�obKd��(���t���̖�OR�v2�t���\^��\N��K��cE�9Zc��.1A#��Uڎ/��D"~��]��ٳ𞓤G��r���������q}�R�Ih�6Zw3���6���q��U#��p�)�on*�̧��Q_/L*�ܩy��;�A�9�wr� �#S�%G�|{��}�]�O�k�#UWʣ�.V/Xs��C�4�\R�EFS���
�_ QIYى]T�j�`;��:��t�NQ�2i������.�cs���� t{���V�H��Z)\* ?Px�a�s6���2��	M:��F[��}a�j(-���(�S��C�"�EŇ���ڰ#�I��v�[��8_J$btH��k!\���р"��
��I}��QZq(T���Cp��H&8r�.MD�uo��tYlk�U_|�87�l�D�u,S���b��{
�g̓������ �X%��©��7[Y�#\�An\}?��Q�ޚ��ak�ƊcED����ƸN�ȳ����͊��ʎ�cg�xS���O�i�9)���K��
��TW	�d�J����.�88)gp�_�'�_[9�gpQ�8r�͙�+���,��Qz/�	`0��]���
���NzwZ!>�R��