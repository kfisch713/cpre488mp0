XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(DL��6����Z��F͍��{��sz4R!ġ�h��NBh.�'}~ʢ�.$jQ������u�j3bt�b������&�Lbi��k����:���quNw`�"�@Z�୑·�M�:DZ��辢N�1���K�8���۟�虫m�'{
�7�l�l&��L�G��:�p���{��e�D��V�W�C���A}	̀;�6q���s,v<s���į�b?���:���LF�Y`�Z}6�Ņ�tֲa%"j�a��G�r���4e9`�*O���'�I:��e�-IDt�������s]�Y���E�db�ҍ���x�H�����p�r��������@�@լ@�}>$Zء-�E��ữd��ґ���e}���ƭ�2�y����$Ga9^o��14�6�iMp���.����nupx$��,x߈����i,��)��2�A�T��j�)?h��p��&��]آ�v��+�{�.Ax�^����m#K�JC��$�4V]����`�Vf^�DZyLY�EoU��(����ݩV���?�b��Hm�� B$m���U�шG!��kw�>�"}o� E>�$|��	T(��-	��=k�Δl�_[�pV��'�ٱ� �4[w��kf��"G}���A~9!ۯ�\j�-Y�f�F�"!��[�x?��=à�0]cJ�&�wq�L�I_�4���LT/���,�f~!�PKEZf����B�Jnd�q�ȥIC�};CDt	Es����VD1�CP��Ha-���-
SXlxVHYEB    95d3    18d0��M�mqkIJ<�N'#$	�t+-!��# ��%����6����NN��"~eV���o�4b�ri�C��q���\����X���m���_�_��Y`��O��F2(\_�2V���p�3LU��v:�\TV����'���D��<q�/�$��M��C�)��	�ӊ�t�0�g$����hE�=��G������1/��Qǌmc&��^�!n9=�,Ǒ�U��0YR����8;� `/`������=��}oC�0��O&�*k-��j5� ���>֗P/���уi,��	�Q�M�D"Su��Q�̥BG�x���s���d��!r��G���A��؝��>*p#f�b��9�@�0vv��+E��й�)7C���7�'a��k|���S��<��sE~m�3��7��vç(u�` ����\�rS"��y�%��-+S�]�X=�xFΓ�Cp�VRn�o$:�R<(���)��sM5Υw]N�h:��;�_���ڱ��"��y�����dI����붑D�qD_��fF��p[��W�������V�5�����ĉ���O��� ��N{�*aAx��iJE6Ʀ�k�$�����/@y:+("t9we�h��s#xv�t�����qo�a�
K�#i����� ���K�E��a��m�P ø���@���캂K֚*�-:�@��Σ֕��U���졾5pq[��]�cL.�;�-}�E�1�P�[��I/��[p�t>j ;w�:���Ÿ�e�m��j؝O���y���˿qYA*u��AH�R~Uxf0��ha�W\�\��?M��+�7%nIW�4�\��^1�i.|�uov�!>M} ^����b`��m$dߩ ��D��3��w:�ccw�U��zԻ
q�i�?�����ihU����w�Hʇ0w�DK��K���d�5���yb�P >>�������'��qXdLS���/�z�7� �*����;��ʷ��4�W>��dHҁ�S8���4Ye�MK�}���B�5�l�w՜��GV��r�i�4����'���L�%�g�~��fM�-3W���l��7P,��P6^���M� ��{ۈ�\t^�2�q孽ߟ�w��S� �Uښ��OTR�Օ{��4��sP?�e:?�Q����'���Ѻ�0Qt��� ��,dZi'Ջ	���O����N �{�G�P�:j�3��Hor@���{o'ow��4�)� R/�J�z�V�2v�D��e.�[���y��jo����Z���,n�Vߟ��!���������ƹ��?��9@Z�yMxK4������]�-��r�O����Stփg���ё^-�3W�r"?����l��@j��W�v/�/oW�!�O�v��a���׺�LA��W�����m!�T=h��H.>�{��y���}��p�W8V;D��h~��t��������O�N�����0䮝 ���D����嶰� �t�ȹ,>���K��m�H.���i�.����_���@��	���%1���s��ǫ���
��ڼ��L�[Ca̓y�=4p��X�[��nk�_ԋ.�K�O�~)L[��=�|��@���~ �8�Ņ�N�6Zu��3���DW)2��O���9Ӈ��"y$�[�0�W�1����D�Zq��P1L���kt�AkC He?i��~䡻���.�pO�<�4�Av�Ku���{�;�N:	�@o���&�N�iTgl.Xg�$�8& "7��E�����������<f�����W,��������_�
cS\ת����oF��i��HZ�et0��/A8M=��V��<&�ہ����#���s�����\��͓���%�����H8�����$;c�C��ę�y�!H���TKw�Vm̆)<��t)ӌ�t.�����kfqJT�+I�n����f}Q�|���Ȗ��J��~O=��	@CAN�8��|֧�xQOj�W�\,Ev��������
uL���c�Hy寍�����K�
ғ������	�Xlk�:X6����~���8��!x�E�*z��(��_�����#�$)&~���Xy���^��ͬ`�	��J\�Bj���-2�uIWz�]A��;ghK.����0�j�����~So��8���B�B�����P��}n��n���LJGqQ��?`�A���v[�%�^���yύ�ylP"rn�o�	�Pdr�[Y��R���$)��g��B��|(H���^,r����A��	��'G��L� �>�vXה�*�N�l	E�D���y�(7X"��C:�����H���W����wEl3?�i���;��?�"������h[�G՗�E���vU��b2�Wu���	�� I�N���ӈ�97��OR����$(4�<L�;�5�f�	:AT�O���7���[��>�<���3�	�6�g�	�Zb���K眉��а�7R�1��yG>����ˏ����Ĉ�h5酢r��W
����7�<w�w'�%�ن����7�憞����dS.�:ʷ�D;W����@%B3�ь!	����L}<��a�ˠ���i8�"�d�6�jjw�.�v)�fK���@Z�<D���B�&�M"�[��%>�F���_�GNA���;����Ҙ�ۛ��9-�p�~
)
s
���P�7o!\%\�hw�0���{�<��H�AX�f�	�j������zM�{S&�܉�/Mܺ[����0�΃�twേl�G^��Ƒ�S�;�r�d����hB

n%ur:��u�߽6~�+���`���s��kh��Oqm�Kk�� ������H#�e/k��Z $Z�x�^ݴ9{�<`R[�g�R��9�K���b���4�#��'�I��������G�϶%��Ϙ��{�:T�l㙬�@$XP_���iE��b^u3x-��9<���(�_��q
�g;ە��x�J�?Z���T
�g�_yc�̀��^\]���;щ�C��϶������\f�HV#ϐOԽ��/@ߝE-<���O��$���p���� ����cnnT����x�,lU��h�"�F�C�
{iP�7��;����Dt���3�ʡ�gg\���0��v��g���_u��jg:�b��l�UT�A��U���s�"����z�>���tZ�YF=�ˈ͘@����jx<T?͍s�:v3�vMb���J5���
�;�w�5��h���&�Ԑt�] ����ò� п�~Ё$��3��;t( �T�Dxe�_j�Ô^e!<���e���;L���/�ة�H@�8'_�(�X����*��M��\�,�&Dt��g���;-;,LIv����u�*J��tՎ˝n���`=S���W�Q�;�T�Mq�X�O�dҨN8w����=�_�� Ah}F~����,��q�K��SwG����y��Ί+NB�1�pĩLԫь�$n^��ܼ�_�8��q�	�n6��6�����2/�{��F�ʖ�;^{ؠhpa�����������6RU������~Z�؀jz\�%�3	>��V!s�NX��)��A�5�by舨��
��OL���,^�y��������MΖ�>/�Qԇ �r�nE�i���"¶Ї�[��m�K�P�@�h���
�y�T��&�~S(쬪rZ����OfX�x��a�#r|E���Q��r�pq$rw!��'���Z��gu��'��H[F��x�U�қ�����uF�I:����8�-�qS���:�mɨ��{d����do�q�HNd1�`��du��������
Rj7�����J��Tn26y���hu��\���Fk蹗s{
h�ڹ�������9`�;�r�u�6����C'1/ٶ��J�/$y��A�f���l�$si\Nt�E��B��@,k�&�=�$y��q�BuV�>���Q���D`� ?�<��+'�bq���6}�m�c�	�POg�?�+��ܵ��>�)��{��;:����.3�8U�v �o{�`~W�2���E>��P�!D5J�U'��hk}A{�a��֦�'e]E�M������0�lڑ����B8>�N��8M*a�:���ͨ��N�i0�_�B���ybȅeN]�B� ��>���ʫn^��z{����:G�UC>�N,mIh©o�
�������\L7�ўp��^0���<79�"i���k�3�f�1_�i�v)�sQhj��+�nA�����ǽ�����ݼ%4j��A���]�k;��+�Q�U2�Y���Ĥm�	]��6E��a�MI0[fq$�O�*klIx���^뙢YSdro�/����gF�/��8ʐwJY�wA�'��!��o�L���Q�{e��]ϙ�"}��2�E��XKT'w�[كg%6�S?�dk�~||�bOd�u��6��O�S��p��z ��V�vI��֟�b�k�F� �w�����GV�5I:E3�,���� �g�؋���_��J�c?�U��=���2�j�`�OI'�������բ��^e���S�.#��.4-��V�a���u�Z�!����B��2�\hK�(;��JM��p|�Z�ꉴ��K:�LD�J�Y���=��l6���2�7�$n.	�e�zz�8��\`;È�����^�_��AF�����uQ��#��C�}j���D���\5������)���/.�XyN�^��H��Fĳc!ö3���mxM���51���Wa���yݱ�c��X#��� zr1��q9�� ��G� R�� �^A��������Ec�g�,|��#'dU��V<��L��kح\7�'�z>�)��󓟹Jա 9��i���)���˴E�z�	�_'6@�����5���#W_jF3uXX��E'��1�m�`�l�S��,�#V�/���%}������z��-M�MĽd�'�t�#�C�5dbW��J�|��� Թ��7�p�w�J�tP��.Q��sk``�a��s��F֊:C������@�ׁ�^��n=�)��O��a�l�&�3�M��鷃���b3͏Z����Z��*��D�-1ɖ6[Y��X��@ó���,Ў�3�񘏃�=ho��kd�S�V�G��K�U����Rs5�>a��y����C޳3A@�瘟w���!(�������������O9�7z�^�<���?rن�;}������u��RfD})�%b큏T��E�r��,9m�6Θ��|�C���c=�Ec2Z��=��S�b�	�eL�����r�W+t���@&�3��VA90��Y��@�-�g0��Q����ar��븴1�Qq�P����y�������~���y�Ԏ��"]B�_�Ճҵ߫d7�=c��p���C!�$����3����"��J������ԋ��MX���e� ��=+1#g�t��m����\�m:����`Pǚ���~��s�ᐹ.6J��v��tG �|�AO������2�%�������r�-t�7�T������8A7GuՇ8��}<?UQ� Sά\g�/����xJ��eT�u@��3�7 ��$��c���"��ێ"���˓6TjO��k�=�I觱��u�4��[D��I#9*i\�bFp}ˢ���ة������ZHxg&`�|6*n�N�a@��]��e�_�[�v��S�	���2��Ҟ�'�N�A~��Ol��L��v��*Si�#s�<�8o�1�?�2�5�j#7�n���+rA�;�e��4�vsS�M?��M�J�q����һ͹�+��9�qi��>~i�j��*@�n?/�n`A�c���!�1�iny�`�闉U�d3���2��34�)�{]X��nd�SD �-CIĸ�c��(�i�	�7w9e�9���9�{@��+ ��6�q��g=���ac��=�������]�)��.��D�s�����T�f�	�R�{����U�GИ=�\���:d^��C��h���m�)Uo�[�Λ ��1i
p�e���Sp���=�8h����\��绯y.wL��H��yݢh�9� q8�*Ls9�>_+��JE�t��'P�V����8O���p{�J"*�d��7�X��d8��Z��N�GP����l}��	]����h�A"��+,s (^�6�HIW&H3Uр�}bU��9�%M-��y��7���^��Y.{0�������)֊Z��,����_��j��5��3�U��f��?JD'oN�7�
��B�#@D�?����B�ʣ��