XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Fݣ6�g5��z#�y��C�q3�*���?eY8d�z>0Bw����2GNLw������9Z��R�>�b6�#?>-��K��`s�t{�g
iE�z*���h����-�O��T�H�X���ֻ�W7��"��ɷ�ug�
^!5�F�;��܀�?��[k�5`�[���-�Ur7����7���Ė���Q���\�ʴ�������&�z�Nͣ��٦�� ��E�O�������m��V�[��'K\s���R���$��
�l�?�g+�TPS�1m.��3q�7mG�o;����(�����/6������}Qx=q�8V)�ȴ��BX���� ��*�ݕ���(���5�B��ӓ'lb�����ev.rkc�����{!�+�5�$0�;˿��b�
��,ޏ�N9(����1���i����0���叩Z[E@r~�(��f��!ۀ�M]���T�S��D��G���Ԏ��C��U�l�d�(V �h�M�0�$^���'�]=���7��&�t萡�B�f,�b��\�t���Ӄ�v������m��fa"oj���GAD�8�H��D�i`�26��e�P�]Q�.��6D^v��Ԟ��ULY�,~3n4�GtnBχ��6U���9����Bj�-�*@͓�҆��TsU��F���'>�i^4��.�18�	�6Z���@�t֡��š�}y �W�z/'��	�˘ɡظ�r�A�1�/��F&�Ar@���Q�p1C��dE�Luz;W�aי��ϩ�2�P�zt�<���OzJ]XlxVHYEB    3b09     f80�S�d���Cƥ!��l���o��'����NdDФ$�2�mlev�W�6|��+��y/����H����τ�⫏Eв<����&���`�{#�/u�.�Σ�ar�wwq��u�PP�e.��-Ҙ[
]#��H��Y���»�O�~��-���S�{���6&?��|�;��0�9��ジI�q�^�(�!�XwC>ϼG�ʉ{-fElR��R���ԕ&K4�*�k'��q�k��$�@d�y�3�AQN��o*cF~�PE���4Z�ӏX~�p�H� [e�Z�&`�J[�O7��*�A�⳱��(�y�x=��Gc�aG&�pUP�@�
�\�Q��NG�H�N�T�溣y|6Gw�%��O���|�8�\w���"n�s�dߎ���n��#�rJ��Ύ�󄱣�,�k�h�i�Џ�$<� yb/(�Zݑ��Y|7�U�
�z����sM��+q-^u�� uiՉ�k%����*����;�XD}��Hp��%=��Rh��OM��V��r<��N!>���.��.��m����m"Q��7'��#�K���y���K�4ꭠk��
y�������T߲�BH��4��F��yW���<�3�H&o�&xQ��"�Uq/�S
��ߟ�妐[�l9D�m�����i�"^�8���JO�A&�L�t���e�!���n師o��!����ƻq0_u�(�l�\xEx��h�4D�qIu�w�im;��&����e9{ś�G�ڻ��ʌ+�D�:^�Zn�^-��~���f�Qf��%�	T�#xqG)��xt�$Th����]`��'�!O�X�*���8��eaq�{��<n�R�(?�t>�#��^�6��|m:��mK�p���Ŏ^h��X��/�I������w���N������! �/�:�i+ !��0����X)J�G+���� :���j��7Y���^��2'T'���D���wl1���Kb4��ʎ�����ǥ������$X.����&63B0�4��Ы4��g6�SUVG3l�ӓ�e��������n������02��-�d+u��@�c�\$������tP)U��&� á������{�D�y��A�Y�U�O&�>�d��� ���&�����=(�yYX�4J~���Ɓ���w�l�������v�݊$���2]����&4�D<j#��ǢE�gD����Ͳ��Y����W��+�p:>Љ4jr�x��}(��gO �89�[�%�N�� Q���?8�	�5M��h��j�~�?���8���% |U�����5� ��K<4_�$�ax}�rT�������狌��a>���p�O�-��q�ڕ�*�������,� ��,���N�T������L3�0�D�mj�<l�N�{�S�Z���7�"��⼁qb�$����1�L�G��R&��?�MKy�+.��C��c�&盪�Q���p���1Ҟw^��П��а���h
-��<b t�6�{�mr���rG����x� &k�o!��%<����Ӂst�=(��x��q�鍑�} �W���Z�,�W3��BdX�Z�����f�ګAw땢ef�%�+�!�����=7ϻO�OO���R�+w��:��\G��+�!��{HU+mw�eRn)�-��Hc��	�z���ޭk_]��N��w�pZO������=�m�ߙqO��7	������7���05 )�n��=��ӯ�1����,�T�M� ~/(���o�U�6ًj�٥F�+�����̜����hD���l��9�^�V�UveE���v<��Q���#�=��=3��L޷���*t��~��0i�և0OD�n��b������e�[�Ģ�������"�\ =	��W
��|s>(ʻ��]��ؘ%V���/"���c�FrBcK�9�!!).5%��3�V%c��|9ճ�/��`N�6�Q��˳:<�K��5�� ��]0t�I��&w������ˈZ�]|mF �!��'XҺ�6�ܫv���U<!��\��������ݸ
���>�3shT*!�y��g9o�?�MⲈiO�U5��{^�/�K�R-hG�&R��f���t !)�9�xS1o�כc�����@]��w�S/-��+9�~ �*ѩ�������Ԥ�����VV0��<������[�㽹�4��|�V�I�+��a�$��i_E
��?��b�!�%@K/<	�e6b�͉�����9[,x�[rշ�"��}��)]*m�1}���� L:�]@��e��:6��z�V��S��UaNg��0"�?՝[�I��Ӵ�A��p-��i<�Z>Ǩ�k��°-�H���q/'x�Υ�XUN1B���TH�X��m5\첲�=`{1m���P;߃tu����:�����~��18It�;I��s�-�b��� sv��o:(-��+~�M�a3��{ֵQ�q��S'�f��[;;��� ��H�-%����qz�[��bb�j�^�(|�J���L��-�#e��IE�=鯊���!�p[O)9�_m�D'�
�9$�K�Y.9��}ՙ�2Ǫ����:��a��'�+��-'Sp�O�W�Э���G���t,(j-�$'�A��1��
��l����%�X%����!�z�J�K����]5 ��%M8��9'�}�~`�����&莟V���T�hcL{vv�E��]�TCU蝅����K7��Td�W���h\UܶJ�=�	�XN�y#����_�Gɍ۸���G�����]����	��L�,z���V�"����"d!�+��.�T���e��Sot/�$ĸ��qK�p%aQU�Y^�o�
CK�B�U:H>mBS�'Q�	�
,M�@��_u�hjBq�U���Ģ|�<�@qmϒ���F&��#肨X�·ق��]�ݚn��^�Z��^Ұ��	>;xj��>�y�q��T���j��jL����4�/�.5�Pn2`�:�,��?k����>ƚ@���r��V9o��o/���FE�==	G
V~7����ц��+�ZB�u�([L�4m��	�非�T=�����up���������b-+*\���|5b���q�)"�=o�W!ė����q���BI�V4giYbK'�2�+c�$wH"g�.�ĎMf2`��t{K��n��m8��}D�H��}@�.���l�}���#�b�Y�=F��4�3=�V"q�w�ɏ�
��턽d�zi�( �ATa�R���7 }lt���ë�<���c��p�	Iƾꃤ�smt�¥�~9�WP��~���=��M���6��{�k����O7?D-p���6��Q�xׁ���ע�4������aj`�W_���'j!Q2�?��vV�]��>:1��Ͻ�m�tNa!
�P���f}y���@����h<�%'�ꩪ��c�.O�A��2�������4V9%��df)$�V�紐m�Z��kd�j�����I�w��oс^�Q�����V��fy�����E�AYr�1}��������I�9O������$l^�E����t�A&A��:6�I�o&�JŶ���[��zy@�`�׈��!���� 0��r���+�2��kn��H�eA����'�9G+�y�NB��3�el�N�|�ML�O�Tz���əM �������Ǭ�V��o���h?�khE#�4���ܿî���Bb�%n��
����L¯� �GZa��'R����q�� ����`d�r�����li��2.���!�x�T��i
����P	���-���E����Md��%Ț�|�'��g�h�מ�F�>5B�'�u	ڐ�د6Y������o��c�nX9�sOk���=��)���'dX�+�/�{6�Ə���v��n�Ƭ[HU�\���ul�d�h�+�Z��)��T��Ң