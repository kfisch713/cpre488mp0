XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0v*���n��T4��T��V�M׆ϧ<�4tn����y6y�F4��u"=t~}�M�[�g2Fp3��:��1�%.
��9jq�&��fDW�Rva�Sb䷽Np�V�^㔳�Ə�b�P.�ke2MϏci�q�>����n�O�T�Pj��l�HN�2NG��	�a#�=�̸c�Z�i�N�����;!FC���垺)�U�W9�Q�i�¢:�­�aL��gcP]sN~���Pr�A�
>���0����.�+���� Rn������� ���g�L//E�8�4yJFTD�����b%����y� d��Ǎ����G�`)}o���.0`�������jw����S�n �M��pXb�'��σw����+����!���K�b�DfSku�pu������tc;H>�R:����Q��R�k���w,���!�������z�W1��QA��6]�3�w<���9L�vI�o�Om�ZBza	�oZ2�I�ݣ�^���(H:��� y�d�A�+ِץz�_�EMmQ���߶8��
Y��J~���J��a�{��%ZO�7��o�	���_#�W�ث�9��0>�'�����\�uXQ[ÔA`��	���L�/���f��d����.�n�p4�����+�����7���ֳ\��]���I�p��ᵓU�
�0Τ��jt�Z���L-by�QU�v��=���L+e��V�)�y�~�{Cv�%�5�����$���.
C�A׼�ѫS�:���j���=��XlxVHYEB    6346    1790i_ �5����H�2��,�� �C;��rkT��ȥg� O�y[�~Z�ۗo��v��ˊ��U��Vʝٌd���g��q�����Cn,���Qo=UH�G�;�]3��;����R-��M�A;��T|pD1�^Ü����f�
 ���M����������c��4i����7xp��ڪ}1|����k���`g$j��z��gS��f;�(��Ñ��Ÿ
�ha�()܄A��U������l�s�\�)��g�dx�Qt= ^%�F�lsC8qT�� �zg*���ڙ�?�H��y��zň)wS�Y�������1FW��;����H��rS6^�"G*�ї�PA*��{�8 �(��YNpʦd&��9�Ro4"#�k֯�)}��By-ϾhQC��s霋�5�7�U�zYz�kR�&�اs��fa8O,m�c�<�L�Q���9���!w�Ũa��F�Ɠ��:�����'d�A�%�gZ�n��ɡ.S,ʢ)�>w�u�)�͢9<��l���4��K"nwOǁ1z�^��в��ߢ��,5���qG�8�^�������J��k�p�^���*])?m�$2��f�}#���ٜ63��_�)�d��H"Y13�Om�D�!_�ѷ�\��\���"IjKL����C0�����G@-�l��ST�>���\��r�����MU-cYk2���ÊT�x=����W]C����h��I��9t�xKb>d��8����0ր`��
"�}$�k�ю��]^�r;@ɶmS��v�drQr�U�ЀK:a��c�־_��-`CUڵ[�W�OM(!B���d����͈/���_pE�)<J�I��s�HY�o��������_c�@b����LsB��kR��K��M��;�k>؅x���G�v(�;HXƋ� ������g�%6Bގ.�d���Bۥ�|�]���ܐ���e��	�U�\��n�� PeQg���C:|�R�b4i^� �5z��ë��)I- A��=?�������e�Z�N"���Rnr�JeE`7�[ ��B�YTN���Nbz-|1<��&�q���O!?��"8��pK8�P���]9ޗl�ֹ���Q�h�v�>i����"Ѱ��wv��=��''�/�sF����g<�#^�.���;�G�I(	W�t5��vUF9��n����_{�z`�e,�
+ .���y_	�˳�)��C &�6�&��-p�)�.���4�y��ө�@S*��x�}駡�IBS���;��k�9Ysd��j�nԂ�M�e?�厈��z	4��W��zү�[��dc�{�L��ʎ�r���N��H�Q����An&��J��ҹ������@�O`����?c���,���:��KH�ؤ↜�6�d�n���H
�JF�������F�;)ꚹ^9S�oq?ִa����#.���	�:��B��6 �r�Ϗ{#I����M�8z�]���H�2T	�Ļ�#�a�vr���I��9�R�h��qc�ld^�:�H�b(�OOC2G!��8wO�� t�qZ��O��	�$/bVei��I�U����o�@��
���c�fwDC�5Id/�{Y֝�֣O!���3��Wa���i)󤇴�0^-��0���H����y	ڮ�&rM:E�M����u�P�N���QӲ��,#�=�d��\n��W��d�տ�axBJϖ��a5/�/���q�i�v�xU&U_�Fh>�D���@w�m�<�#����F_yZؾA@zJ�S"8$���F{����ك37Z��R�������t϶���9j�:�QM�9�9=��q����'��&C����x>������t�D4�&#��mdw��Ɲ�k��P�<�U�B}vRQ�AC�����q?��P|�2�7+��V=�ѡ1�t/�>����b�r�_�ƏY<+g�e?1���y�'rxF:�sm�ϡl��q��á�-T��v*��C
g���g��x�}~�}/Rӂ��0Yb~w�f5���_P�/D ���r�p�����Px���ڳR��tx]�������^RO������7�� j���p�b���8ʒ���d���TԱ����� ȶ����V,�	ˋ<y�2���AR<(��QTVN���2Ob���|Mk�/[Ԭ��3g����y",�哎�H�wz�6�2���Z�1��\�����a����ʙ�NAu���L(�����b���7|��Y��ƞET��esc�#�m����:[P����&l����K7H�w#��v�k�Oz%�L�)��7��Aɫg�kk4�;t�Q�j|�'ߏ��`�U�cF�r�T��R�V���
�bHI: 
��kօ��؁��M��/����]�%��kE��s�3�Iȼ��v!���Z	�>Pr����m�4b��'�`
�Ü�K��?cB2CAɸ3&}uס0�t���`��� ����cm&{]�y�'���!���7�|,���Y!:�h4_���×	I����-�\�SK��2��~7Va]�@����9�m����\~�!�.��E����-����߯�;8,�,�b)w����866�1�*�(�7���&
Ҽe�����v��v�P$\���{�J���t�+Z&�r%c&��Ā"4^���? І�U�:q˙�	t@J9�����[�*�Q6���e�(��������K��"��{�k���`^�ެ��6�[3C��f+����+��9y�#�Ű��OwfW�w���R�.+�F�Nѣ6'��D�T|]�?���~�Q8��خ�5�PN��^N3���Fj.��=��ٙ��	�M7D�KH�.z�D�픹�wOA�4�R?��ހ��NB~�m�暿49qMS�,�bwe�{؉F�cm�{b���z'xܨ�R/H5��#�(���e�;w�B�F��2��2� `�K�f�8�R��;5����������2�@4]л�V�8������V��
9Y�X2\���2����t�Zc�I����De�����C�.�.$�܉�f�x��?�!%x�ti��8���̩&�w�r��oA��v	Yh��Y����Wp��&����{�P� {�[ ek���]B}M>�5Qc���O`
�z� ��FN����zM�5���6~�$�5ɰI�-����Uh��*�T��0}���)�$b`�+��.����3 Ǐ���+	���U�����fXx��Y�9ٚ��s�z+��2�ѵ�b)�
����.��Q(�֮�B#�P���7(Wi�W?~xŧe��o��0����5QL���;�h;!���J�O'a"`b�RzQz��B[�O�`��Bk�幋��`�}�xTa�r3����0L��w�����IqoD��3����{a- ��T�uW��0&��'|_ʼ⭾�BP.p�5F|04������16���W�?������č=����m��w~w�!�
�(@rnt�\PVj\I�"aQg!�]̻��~�I��<�Wl�	�cE��B�W�ӽs87:�2�Ei݀���JC����dв�w9W1x
���g�+��őpg	���h�/{M�Z����������08�tG�N61���y��QJ��‌��Ϡ��11��y�Q9A!�*�`��mψ���u�&�ɯ�D�d栎kZw��u����SH��YҜ��"'�}����f�:Q�yBѳb�2㰸�/���?����b�Ct�FN�{fE�+�6_L�cgݾ��q$��p��S?�+�&%cW��΃\��Q'XnU���,��ec�s丙��w���,T2��1/��u����6x����?�9嗌�=����;����"+��an=/��_���E$&-�����M
�=+�{ui<K��;,\�N���`�ѩu����&ű��&��/YK={���f���
%�b�=x=u]��v�ϐ.��݅�.�ܒ�R�L@%�6x&+��`�MW�+~Ŷ��q��,�V��PZ �ߞ^Zk��Q��mm�U�lMS���i�!<���o��_�őȸh��^n&�>s֬g�;s(�A�����Q&�I�Ѿլ���{�q���F��@�5L��)]�����5К��+��KI�{ٞ8F6i�=jg@O���H�a#j�nx��N���c���S�����(�����U�G/�=�����[��ao�is�f��r�C�t��Bfb-���s��	ϡJ'?O� E؄Ȕd}��E}FN��G��h�T�Z�W��}�?�j�v����:�r��F@O?lLp���A����i���{�ډ+ۄ8S������O�|�����n�N��RR���ڪ�22�Ʊ�xA/�e<�5Mww�E���p�m��*On~��bTG�w�L�߽�6����j��xΘ��9,����gj�rO+6�[�,�ߘiB<g�5ʟK�5+��f�!̒�6XܨX6 7����P^v<2d�t��n��-ފb ��Ā�|z0�o7���3�N���=kUZ�~�B��B�iPU��M/=l�!UǕlB�
�O1��W�7r����� �a+�i��d���.�tI�L"�6����?�-�Y u�-�ӹ��JnY��=hD ���_��r@�{wD˪m���� 6����j�PIեl�#b硉�.Q���aӥ	�]�:ŘV�DQ��Ek��s!�%j#���_`�A����49ŕ�ѳ$�`r	�٩oVz�h����4�uMy �q�e�����
-��D�o�eq뽗�\aF��/�D!$|�� �ƒ�s���^�h�^�x��p&��r�(��_r*<�^�!j��p�����$	�R�=�pL�b� Ռ�������~CK6)��f�-dwf�.u�	�H@��ahG���l,X��2 �Ч)m�������	��������� �c�C�|z�A�3�7G#�eXVC�/���azz&0dW��d?RP:gbФ�������U)�{�[��b0��Q�Ro����s�3`��Z;�U ҁ�knh�~�˱e�ov޼�iT�{��qk�PƂ~H5�k�I+�;0�D]�T��,�v5[ZY算 ��������4J��low�;e`�`2*�*���,3(��߮T����D�F�\Z:��%�<�]�	(85�r-<�72�Rj;����Z�2M�����@����v���S�7�����/HS�R���Z+S�2�eKU�~>��}��0�:�����-�����,�D,d��S�-wRR҆
��{{$�v��J�uɐ��$��M<�)b�����v+�쬵rV���kv�q*$���R��Q�a���Ǡ���Kϗ'��I0�`�z�4_6�m���� �N����X��.�U�	}H�0���l�
;D�� qm�
���j�D;"߃�
�9Ŀ]~���"ar����υ/6��y�(�=��EC�����u�ѩ6-L��C�I!���騁s�a���3䒪lO;�.c�E���H�J|���Y��_�ØÚ`�1~��7��j����v���B��>��җ��??���M)U�T�,�M�M�1ro=B�c'c���jh.�q	�a�����.��}pd��y�>�*�z֦��!�8(�`�\��AKe�*�3_��$� �u����pNyh.���1�t,d�:Q.�#�R��nlv�O��F&�� 1�'��-�x����O�#q�8a>~�?�������SJ�[�� ���=C_@#9�D%�|\i��<�����֜�+��d�0R*	��} o�Cɇ��Jo��� ��CQN���]5j��O�cK����&�c����*��e�2��X�t+(G�C��0��Ϙ_�lz�q]ę��v��=�=�Ę˃_������wt�׍��qjF/�N��Y�l"ђ��8��-9�t�`?