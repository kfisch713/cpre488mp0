XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Sf���3zX#v���>�.���o�Ȉ�e9v��0JT��X�ނz(S+*Q�7��]���o:�|�-�C���>m򡜈��f��/:Bm曨�i@t��_����/Gsg; �<C�노��x}�3ݞ�5�E������uN����@�@,QSΤ�U(��T��1D���d�V�����Y�d_�n+ͪ������最��]�i��GN����]��`!u���U;	d�G`��oVQ���63x��8�y�Y���1I���g�q��G8!.�Z���GwMn���:ȿt���?C�:G�U��:n����`�� �����S�%uؿ���n�����,.�Xǽ�v[��[Q8��Tb�1f���S�&��kgNud�����XX��Z���쿪��:�B�r������:,��_/�̤��j�o�o3�x�܊U��N�7�^'��3D��Fѻ��+��j�<z�^�a�����T�.��@�:RRĝ��Z�(�q-��J� �$6��|��käԷ�	�D�t6�] ̵2R�\bLf����Q��_�����|@CS>Al��.v�ޘ]�Y<{�3��,yAF�������H���̸|5��K-�j�H�t$�ɟ:�=�T�HX���w���tV�I$�D�$��ҵ���u�ڇԚ�sN�G׵���K�.Ӛ�lk�v1d�<�;��ā9���c�P��wW���i�b�.�4�'�v�PP���� ��o7�>�}_���2{m�^6��CGXlxVHYEB     f6d     6f0��M�ֶ:�тW�]����9���!
Hsh7�:5��CW*=���yN-OT�,$��/<c�r���yR��a7��M)T�e^�{�dѦ�q����Ѻ��j�M����t�x���įc���Q������8#���$�TR`r��m�#�r����Ö�F��R{��ќ��,I��^�h���?|�r}`�zi�&���WFmG�bM�ܑFV�c��Y#�L���'�Fa/+���4�^�7}C� ��nw�|ŵ�4�jE�q؆�`�}��,���1c��_-'r�F�/cݼ.c������s4%=#��d�J�,5ᡈ�D�yX��}�h���}�&۴E�/1�uğjdJn�p=$I2F;�a��4"��Y��HF��b���~�"&��TgD����V\8�!��k:�����F��>���")��d�0.�-f�8
���B��9��~xkd$ݮ�Gx��I5� 쮥B���@����O)ѳM������/D1����'0u���ߊ؜�o�����^�pЧ��^ݼcL�ߌ�RlLC���^�,G3�v�`���B�(�M��U}�1�U3p��~s�#�>�@#��w�Ѵ�$D6�S��[e�L��F��(_Mqr�Ԇ�Zfd�˻G�1��,-�hj�0q�W�(���g6	_V6okҧ����A0�KMѣ�֗X��=�BWԗ�M�F�{�����u�1�*�K����A�r|4ُt��S���y��#\�0S؏�G���)�g�,�9�r���q1�j�*6?&9v���>g�N馦��*�E�?�F����2Q�q�]�)L8J-�V����������.�[��$n���qq��A�L�M��<���Խ�9��J�|j<'�o�f���=��q�pCӬ-:���2���LS�M�Ӂ�'�$�q�v�1����|\w@*?i��24��=�*aH �f� ~��"�o�R�	`v�r��	>&PW����T^������ڒ���<�@�@ł�,�yաO%Y�"�%�[r�C?�(.-/>�ů2��E1ߨ|u��WTL�nA+O�.�!�;1�U�E����3�+�c�A�a���f>¬�/�����:�7�=M�ʶT�xg旌�|.����U4�Ci��
j��2����d�G���D<����,{���?y�d��YC�S�� ��yw�;����?���r��?�N���{���� 5�N���
�!^����i����cy D�}���U !�]Tɨϓ�ziE~�v
�&�,���ǟ��9P.�¾����Hi!���e�"�]�K)��D�x�?P���G���L�(1����	V�Y�'���8��Hˉ?b���ӇC�3����娌�UТ�F\��Q����Thic����m�@1]�����xn�O�n�Y��<���$A9(]�5Nx���D�\������N�h1���f��z2���]8=��#V��^�0��t%��c�F�2x���HM^�}'�..����= nW�"�~�c��!�؂���W�<	9^�3�"Te���4U�()%>ǃ�p� Q��&�s�A6��&����a���k�/2f����	��S�z��n(��W�J�h$���~,	x��lJAu����t�z�Op��?��,���l���y,)d���*ΤqL/����r_�h�]��ͳ����0Z��>��#S�&5n�'e��x���..�!x��Y"Bm����M2��uA�)6*�