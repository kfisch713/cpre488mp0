XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���4�Ye��h�-��e�z�{�p z�Ջb4�0p	Ic0W_�+��a�$�)m��a��n�Q���2�pR�I�'k������Ji�Yh6bU�ˀ!��������1�̆*dߏ�*u
#�3�8}���Fq�U�]�tŀ����Ƅ���3���轪���I��_6�M9p9"�{��P�-kY� )��h�xɃ��#��j�hǭ<��tPo�1am�+36I���n?ٜ��$�V�?+C���=��'�ߝ�|����Z8-�2�f�76hŉ ʊ���=r���M�D������Kl�5��|��w��X_pSܹ����E�n��IO*�͕M!�_��"���d��F�z{��/��P�����*v@�ۀ��Վ�ִo[������ဢ]4�@�d���X��Ge\��~�E�H��\<VcN���������*��F��;�Q�]�Y�x:K�Q��q�F���0�hA8�_��.���H���&|�9�Þ9Y(���	���$����(_�h�H�}g�'����D4���$)e>�s���é���ZW���J��_r����Κ�F�����3*y���*s9�G�|v���18�q7r��$h��3U���/��8Cג�oD������T��rEpP^'�g�y��
#8��C�^[i]�P�F0���;�'����T�V*���{��BaJPJ��p�V@�EP�oF?��⸮Y��,�^Y�IN0���ˬ颾x�=�������XlxVHYEB     f6d     6f0,�a*�tƖG1��@����Ĉ�2�u@~��*�b<?T����μM����:�4�IK��>�Рa�c�^	D;���΢?v����e�7���_y�2�����6�E����:�c �[+�5Co�p��X�}�
Dq�%���c4�?њ�Q�(�����9�=Ĺ{�aO֠�Rf������\sk17�r�ɧ����Q��C�+��aS��#'"O��Jd�/��񓄠R@C�̛���Nw��x��ΏTq��=�+����������t��� 3NĒ�z������+�"�`E��$�ׅ%��q�g��V{!ˀ?��r�\�����ċLI�#�Ү�g�`����sZ�o�C�w��gt�s$M�zN���w
^@��mUQ�@�m����@.n�a����qJ;⚃ELa�qǹ=f�Xf~�䘂s�����H�VLō�d�]��C���1Z�F�O�>���z�J�b���v�x����d�7�M�On�iMXU���(-:y����}+��;(��읛'�֕W��XP�
�H>�v9aY�~�Q��qY�ׁ��[<u�e�œ��ܢ�Cu��c�cV`n��y)��zG�Ն�4�a�NT�F�c8�/��"���G��)�ήsI�R裇���j,��s�&��9�ӧ��;m�Ë-ΫX��-�����tPۅ���m���s�[�o�Y����=�w���:���{$rm:@Aء��+Fb\0������g(!S��uϳ��@U�?�����72}Y�B �-���&�h�/Yn��Dj(6����ڌ�lߝ	.ߋn�I�(mQ]B� p�5��� \S���ET�pR5q�~�[I,ô(����>n�M9CJ�\"���M��^�A���?�k��L��@c�̒�|�k��H�3Z��F	q�F���*�Q���_n��J�P��Ks��*���-���-︧ ��g�$k�M�}�"Z��dU�=5>���YO�*P���2�eHm�0�pD�o4*�s��S��z�S���3��8Y%N�d�9�V�D��_P�Wd,7��c��k@@�
*��Sâ�9-�}C�R��Y���m^Q��!5�4�`��޳U�{���� ]�^���Z���i|����+䜳<��O���lU����G�+SH�����-xIS�MV�h�����T�:(:,���[��x7���\��e7�#�:M'��!��i
�n��ab1F���Xz��$1 �����5zR뇛��Cj�9����n7A�c���wɊw&�D�-���Yȡ�8%��.5��M�}����ы���2<|@Z� �ɝP�s���E���%�ё�d�ށ�ub����>��q��Hz~�QC��ׅ�Xݝ������r�G%$�� �-��m�`L�o����l\v�Y���jQM�����po�>���&�j�M<{k�i�E�GP����:��ϕ�,���u���n���.z���%p~W�6W�,�}�`AI��Q��o�-�2��a�_F�8G��B�f��q���'J�t�߬đE��-���@�����=����c{L�Ot���H�j����ɹ�n����@g�T�ԛ�/���ٺe����`xa�����G�IĪ�u��ւ[��Pl��*���8�`SLf3��ȪL��В�ӕ�����tR=)�:6��8\({�ف�(��#�L�LS��\���w��s�k7���d�2��b/��A�l�6��