XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Բ����B�$v��̒���񧬓��_�!���8�w�Ƭ�Զ�-� ��i�q�O�����(ؘ&��A�
}���E+�;�]m!�67�y�v�HԆNw��v@�y���87^��·D��� i6�H�n%ظ]���ʲ[��3|,y�Tކ�
���MV�O� ���&ia��g��@[�>��(R��ja�%,L�B �?/;�IN�5�Β�f�L�+�-�X�y� �V�"d�6��a�.�m*��-YD�X�`��\c��|�d�N��7.�L_6_���K�Z���;���ΰ���
C>2�'|��U�yȧ�]�i�_�޴e@�����
4�9��f�0��@p��L�	|u1̯�v���v���[�gbb�^�SV�K#�k炸�����Nͺ�G���m̎��^�:Wh����\�O��=Pc��8|�8yt�|�W�����Zߑ�����_��*r6*�l���j�E;��\�Gx����C[���=XT�k��zV������Ƞb�y�&i.�bKP���c��C���[N6��*��5rAqM��.�-4�V�՝kO�V%���8��Ƿ�[W���f�m`�Ф[꤆�+��gY(\����c���z%Eކ/y�n��z;�xR�ecmW*f���]S5r yߕT2$�+Y(�hX�hv�!碙���6��RK9]�b�Y*�W��و-����۬YeE>i��� �d���*�P�ӽ����6�Ti���w"����%���KXlxVHYEB    3b09     f80�$/T7������f�EJ=���p��)�o���LK?����~�>�����S�T�������+�q6������\&���ҼpF������6n������:#��f�gu��Xi=��9�!��X����ڛ�� �UZ����}�1��_nX����L6�,�Rg��n?��Gu��r�
:��������Qb����G�����|�a��2vFn��?TSr�(�a��5t̌����)�#�|�q�%�s�b�ZH$�T��x(�XJcl�0��4l���!2jC�� �l��;WS��F��>�fƣn��o��?m�M�'���$A�q�� ��֕k�ն�kbp�Z*��r�֢�)���g�8 Z�� �ji�m|^U̽��C�{@O���ܟ�O��Ѷ<wDI�+��l�H�\�{�z�D��Y�FM�X��m��gi��Z�#;�"�wiqP�'c�4Jc��M�+��������BՉĲjT��Չ#�q��Uיm�4@(��b}kw�^���+��P�r��3ʪ��{ d�a�~�0@�3�Px ���O��V���l�rK&�ײbD��������$�y(�4���Hy�j{��������ᱳRj����7{�k�.��`����"������{$!��M�];]��Y�ԿP��1��d^�����D���ْ�`"M�����(��`8�9{��pۤ�2g��n���A�`mQ>;���Ysz�ME�E�R�P5��.9�k(�4):�ƾ�1�H5����D�|��HC��_9z45w��� ����>��xPu˹���h��WR�C
	�����4q#��k!&tQ�)��sd��~t_͛��C�.�������t�������f6L�,0�ٚ�	�5��M3��ᯨ�����^壘5���2����N�ZO�|h��7�Tk�&�db�$3\.�s������KQky�.թ'[�{�S0�(�g��y���s�R��ܛJ-J�̶��uF��$'o������G��؛	����m���+����'))@��;��3�Of#}Yl�B��Ǽ����u��k	J���b�����nY�f_j��Li ��[!ݛy�A�2Ѹ7�������w��l '���� ��p���3���Nѹp��I����s�Њ)$y�omL�}�K����"����PMH�ub����t�\O��D)�9���%��� ��p79`�#(�0��=��M׈7B���Ř�s��D�^}�޷w҄�(�Bc�T��tU~�YE�ı������dG��ѱ��xf��`��1a��~i�:�c�>/�Z�`�w秡���7��I��3L_�W+�D1��[ A 'u�Ҥ^0<E�V�#ej�G�>�@!|�0�������?���f�ʷ<Z������W��>l͐�Jׄؔ��*��"_�\����2���{��գ����j4�ƥlՎ�����>M�'i Z^Ux���Z+?�r��8���B�T`�b\m��.�X��#���i�?���Ly���CV�Ye���:�\�ZK>W�|,�8B��fV��i������}�u_´��3����{Y��O�Ye%����'����/����w�֘#���[�xҞ����V�PU�0���}ML+�u�������<�Y�'��r��|�bU~ck�y��I1�]^P����5E.Q|tm�|�o�	�(��K�d��{��M�X���L�PܨA�@}�[�6dAkI��>sz���h��R��~�0q�RS��&�6�+�F����`m���l:	�"�|����R�G_��Jb�Ku�w�"�m��`�h5覘��48�˴28=�KvbХ#,|��̬8o��Hoh�8����Ɲ'(*�TH�����y9��JÊ,����ߗBW���y�G'n�d���(��0Z�~�~) ňXɴ��[�37�I�#sv'��g.. ���NG���]��2�E@��e����*���޻��	��ڸT<X�ۦT��"��Ew+��������aF��Oh�{��=A<��`�i.~U�e^��&����ۍ}[�m� �0Nc���N�jW0#��V)ps�}n�u�X��"+$��q�o0��^I@��-�y����>��Z�g��K`K�V^�?lPa1�"]���C��d��b�������d��v2[�r�@9��H�����D���}�_�z�S;��ܮ��i���-�[Q�Aa�un"R����ךK��V-�
)n��*�����*�M��3}6H�B���(Y�+
+\���"���RaXĪ�����%`4ot,����6RZ�$�]nƺl#�D���,��7�|d�«�PqD��  ��3Y{ Q$�h�%�iú�,ˀE~jKqڈ���

KH8��CW��%D��8�l�����69�~��s9�
�d���$�1$׆���nHq<x��;�H[�l藭���;lpe��ء����ʑ���}ؕq�S��_�3��'	����(0����K�kF�S%�8)2�ɠ��;9�h5V��f�aŖ���TU�.��d:q�
�nU�k���k�Я:h	{�����TT:�Q��5%F>��N��y<�Z}bW�&��v��_M��f���	�Oв*jjH�b`,�A,<,NS�z�0~?���V��6֜�>&$�I���3�6J0��R4n^���"08�L��8�YC�ڏ��0�;����~a֌�Pj��(��B�t|�o�*oFB�Vh��q��4"Ub����g�eʑ	�uL�Ҋ�Vfذ����M��c�y�{� (�U+b��2�%�#�CYQ�ɠ�2�C:5	�n�?�(��	r�:����Z�#%�͙$XA��N�׋\r�;���$��U�5��ƿ�����ܖx�y���t�D6�����a�m�B�G�4-��3FW�%ʠ��[�_�Hw<l' �<S� {�w�4N�zp��Oi͛�*[�(2vlI��a�
MT�;��'�?�u�f4�m����2�(�t�r�I��P��;u�����]U'��"Dpfǰ�*���ehz��;F���)E���O���Ҽ$v��]n���4p��&���׶��6��8C�bEO�g�u0V)ž���[G���-�Z&��zI��͏�eI,:�~wpU��xm�R��'���YY&�x[����zt��&�w����F�j��D��p�����m���h�{gZK��[�};�= ���@�5b$v@QbF�m��*�k���j�Ư�:ٻ�j8��	n7k�JM�����s��s�C��`fek�̒g�i�����;h)�m��HD�kvKr�7,�17|G�]�A`���:b��;��G���0lb�	`��~n�Iv`����J������olI�K��,��f���?U����V�0鰼i[�҃���I�<�`�sB���������;S�܅����]�^
��:.b���LG�D�+��V�z���s�sI�o����k����W_�s��̕%�T�B�:�<..�<x@uTI	p��K'�!H��N���:��&J�0��ғ����0��B���F�~qm�۰{���/(����m���������)��/
_��@���f�Hj�c�\��X�Э���r'��> QX�_$6�$:/Hj�ī#Ū�u��tY��\��X����&<�8y0�#�m�D½m�޹������E~vё�����c�Ðb5��2���1�G��S�:E���e�p;����
~\2��8�L ���l��}Q/�g ɢ�2�z񹈈tə�sHk6���J�jj�/����eo:���Hո�|lI�[��#���N��=�w"�3=�ģj�A��ݒ�6l��S9\te6"}H��ŮU٣�+���������Qv�LT�u�
u	��s���