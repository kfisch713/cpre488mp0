XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��BnWG�c�0z �?�Jٺh���x5�]�yM�� ��Ǩ�i��J���LJaș���U����]�$V�@!S���`]��3m�r��F���E0c0��!�h�o���zHI�jl��\�q0��OD(Q�����*`���v���}�k����'���d]V�b��.K�AOt�!����!q�"���]���[��fF�TB_�7��� U�䟁u8��=$�E��}^�U)��6L��M��Y>����)Q�B[C��(��V��I�	��q]��UyF�<�����0����^�W�lD����I�	]C��'�.�)�r�m�e�W�P��Ʋ����X�c���i�ΫV�E���'*f�ǟ����V�?}�}-BC���`*��\�����D�j��[[әd�����0�9�)��4��PF$�bZ�Wu�=��ɟה�9�/����K:)W`�y�Z��R�-��?3#�@�"Z�V?�Fv���+��K���o&�֙ %�"p4@�O����_i~>��!7��-���/dhL�ެ<�)��H��I��";�g��iMC-�t{� |W�*��u�P@h�m�'����أ�~լBP��\-FV6�ɱP����)��1<��l�F~��g()^J�e����å����`��^��^��q���hJ-��=��(>�'�#�)�Ù�1d��ۀ�3TZO�&�<Ɛ���C ��b����x���``�/t=������0�,�6������U~�+�h�V�XlxVHYEB    b3c6    25b0Fy�O�S<���Hy��Q��T��Df._���]L�uc��%��X�k�_*�E�5�'��F�Xsiڬ�$�;�(��,��R����JN݌���� �������z����hm� 4p)s�C1��ܸ#�U��2�Ɣ1M�]8M(X���C\߀��.�5Qkwu!��Et���\W�� �y���j��J��uF�
�BvN�6ӓ\�����]'�:�ӹ�>)�[u�5\���й���Tu#�"�Y�dA�S���N�6��<k'��H�G���S���̋�oO	�bNȪ��/�<^�MOG�.�7���pG�8������p2l�,�B��x��&|��eԡ�T�2=�$b�e��Y�飳��4ܻ6xvʁs�\"�JX0r�}A�Sp����?�Q=��Y�#��H�(
C/��B��=oG'- ��O���k�i7?���|��M��A�7���Fz�Z�i��^��a���f�s@�H���
3��.i1�#����J��R3�<c*-`ReM��׭J�=4�M��#@��|�ZN��in��j��u9��K���:���.� �y��#T�Qx��ҁ
PP��O��BKn����ɷ.!�c� L�I��T�B�ժ8Y������]̗Y�yŝ�g�#�(�~*�W)�G�Tm)���)$
�����$��7?IN�-��e=y^��52G�dVQ�X�3�*n����Ij0�1��%������F�)������v�To����{��DF���*����3�u�1m{�|�0��lI�aE9�	��|x1)$�[Q�]27'�tM������lE^�?�z�-�`�ɌE��ga��z^�����&:wR���F�f�>q��Y�LL��m` @o������ȭ��[�s�\�������:&`��S�1��6��G�7�W]7�WHcU��#�e��얠��@�?������0+����>�U��������yt�[���IJ�l�v�
�^w<m0��7��_:��^|�L��ƈR��)/�҄�Ԛ�Z�K���QRp���}��A$B��_d*/Lf��[�(e�-\A)�
�NWF�>a<FV9H^�j8���~Yְ�A8<ݝ-��a�����% ���qO����T��9 ��c-��z����`��n/��L.h�O�^�4|�oN�=��*
�3�(�۲��A�J(�ߧ�;�ͬH])�q(��T�r��)F�
�|f�����Mդ8t$n�&A�`f�r�ݵչ��ao����er6N���byXL�`o��C��ҦR�-8Ҷ��>�@�=۪�GQ�~�{�֘�Kv��H1,�|S��:��Y0w�t���/j��T�-R���I�����ي�/��>�h�6�!B�V{>рD�Q
��1�^�ҖG}����av���.Wa�rU�ǃ��M��75<�q�f6�K��mZ��T۸�vE��HN^�^�CT����@�q���ϕ�V.�]��s&�\{rqT�E��@�p,�Ձ�V;�����Y�������6���'����63T<Hu�����Qoq��}�f��s0"��<��N!d�{���϶����v}l����Qm &-��Vy�3#�	�ۉ�w��b�V����G*�?A^G��;�b;}��������H�H��Ya	|	:���퐘bQ�tC�n)b��݉I��$#^����7O���� S�ά慒}���E��V�,���e��[�����!hi;{:��/ӫD��ܐ`<&��7��+bqʲ�1���F&fy��*{W)Ǖ���Z�*��)����9�ٜ�/��Wt�J(�K>q�?�5B�orR���,�Zc$.�_p�إ�HX?l��W�z�Nv�ˤ����(L1��ޤ�����/�����b@0#�xÐ�	�cB�e֚%��o�=��=�����rj�������)�1m`I+D	d}�+�����v!��:.��¢��U�l��{����+&��c��,�G��>���8��M_N� �ބA���x�ՙ�ZvU�]+ѕ@,�#�V.���|z}��ȕ�dmV @%&
���=2�?��̛`�af��K>6/]�rc������w�<���^��O����"I(7�o�t��7�Ʒ���3H�C�v8%��3Z)2vX�QK��s����-[�ҍ����D��?�5��P�4�+S�s�����tV��^�'eޠ�!�,߀�rk��@��2l{�5�ý>�&�Q��N&�����1�j�S����*�=�����S���=.ږ��>��V�����ei����
-���_��<�v�(S���e8���qVlm;솎J�ۀ��mE�li��K���	�)z
�F����9�1��|���M�Af���{�ן���`sD:̔
#�v�ݸ�"���t���L2]|���{�2vJ�� �#�x=<�Őr��G�0�L3DUT*�O��<�^J�-�~Ȳ>�6����)�C�?�vI�H�j��P�0JW="�ع�ҵR�g��*���y}R��#y#U�a ��������P���
-'Lf!��s�l��%kC��Ʃ�<$B�?Y�=PZ�e�G�֮$��K���O���ڲ��A�7Ӱ*�I\��#/��!nM��Mmv��4�U��rYMn�ۆ&���@E+ܢͣ�%�%Ov���
t����k뤤�*i�X��K�/M<���*R�n,S�ǌy��8�:�P��;w^��T!�=�Zk*��<�@����V��SA]�A�H����o�ʒ�Y��!P���c��ܞ���A�?�9���){T��&��Z1v��jww���{6Nk�L�5�a�d�N���AP�p K�k�l�bّ.�{?R�ä����g(������ul!v�g I�|6�)����>b
3��*����jD�y��<�b�[���7:�v�<S��!^$ִ�3��lE�:,PM�����n/d߸����ۑ�e�p�I�c�}����ʹtb�ej�%�{rƧ���<i���(ZC?�?�(>�m.��k6{�D�Կ��y�`���Ƚ�8�t�����rD�o@-`keN����$�&{�gy�'��]F���&���ozu?3�3`[Y��܃��'���*.���sfF�+�{ti-�i�,��E��s��I�}C�ׅ7T��ω-�R�ߙ�۬<]j�e���>'L(:�t=�b�dMF�fZ#���ڇ]�{s<��28F��`Ǣ�>�\A��[����-�R�ը^�L�	�YI����Um0�V enurg��^H� 
q�%�8Q�i�0�����-\S�4m#l��������ӡ�5Q[ލ��[�G�ZZB�'�q+�R�]@������$�Y�,f#8��)a=�'�V�~�yn�����K��� �:�̔���C��M�����t�=n\�M$�W'��V�{`ɨ�ͨ�b۬��F��V��>.�6L%�sn�-�������_!�wyȶ�LG�ki�H��ӾŗK1r�Y�yX�B�+V�0�#��7��0����C�:�)��S�u}#���`��@q��S�
Dr�beG�D�lCʤ���c^F�L��ԚS�іx��-5���+5A�ś��L΃�g{jP'u�?��ۅ���N���NSrf��
�֔�"��3���n0X��9%|��߅�R����N	�[��!t�"�v&vy�'�()�Čt�V Bs��>���c�<�3	��f���dc`N��OV懂°��ދ���:�9�Q��E�bF�F-o8��������c�<��q�� n"j���DQ��yzO6��5Sރ���`�R�!H� �������F�̈̈́����n�4��4���$������	Xj߭ח�f��px�hP
�L��)�]*�Z���`d�Z6��3���Q\K߿���ⱑhQ3I��w�͏�-�W�UF�J�����[��A}�?���w��T���̚p���퉅e/�v(͢+�Y�XG�ִ`K�u�����zr YII%�����sn艃���%��P�>a� ������"�Gj��r�L��@u�/��;JL�h�8��cA'vd����(uL;ș�z��
��-sϜ>��W?LD���rW�O�JP�C����r8�Y��'>�һ��>���Ώ
�u!�U�,
�O��ܫ��u��%�銬1�k��]�tp���F~uT_�*"d�47aQ���0O����1s]ث����	�\=9p�aG��L�#��I�ܭ�
'T�(\3�W֣�«h<�JT�+AL`Q�߿3-�j.�ڞ��L$)@���9J� �5j��1#7���b_YA8�C�.]ßM�5���M7�u6j��MV
���A7����6(����UM�>! V�V�9o�,�����7��2~�ƃ唷�I����a�PМ�c��3q�)s[�Ќ��Ɨ��G�E�T�`��f�
��(�~V�ĀOz�4%@���e��*I�l��#SdC �����1��a����U�,G�t��!0y(�.���4ogG<�J���9��,42@C�Q�������Yz� ��D��n-�,�,K�}jQe�o�ϝ�z^��ODa^=�R2�AKU]�k����x:�������Lգݙ���t������U~�����a(qS�g�����k���pcW�� �G���B%���������pVʛ۔sr9���Z���Lo���!p��w�V� #�~<�۽���۝G�ACB�}�~܇ӖT��D^���^z�f�˨��٤=�3���n�C��� �F�[d�Ω�k ~*��x�ǃ���K:RE�����֦=G%�����g]�u��҈�+�	����!#h\$��H��DA�J�Þ�&������*�:�G�3��qb[�䎚�(�k��!l��u1����P�oA����/+�,�g%�a���+��F�5�&��U'Ay�Ge��B��O�l�Y}�E�ߐjm��t�Ud��\_ԓB����7�j�֋��Z:r����r
(�WT���IV����� �����u�6(�J�|pQ��
�XV��-�#۷�?��i2���&e��[RO��=�yr��PF�܃��h&/�E�&��*tr� ²I��+'��zg�-��{m ���SQ���0�mL^�4��A�d8�;�xKj����y���!-�Â��]���<�壑�Ka<A�������1�R��Y�>M��i(�2��y��ĳ��ũa��e7-̪&����qm�lS}�]�WX�(ѕ��ܢl�.!�A����3���4[!bj9��P��\g�G9�����߆��^�!��y�O�c���+�X%���6<<L�P�ͥ���(r�i�s����r�3�w!���$�� qn
2����C����I�rE׭�/ <��W���<��_>�80;ݥV�`g�i��_Ԉ*L��Yu����3�($ul�qNh�`���q�˱�(����F�"z�rhy�D�5Ŏ�����~����]�ڟ�c���M�j���贰8���DA�r�7�Fݦ�L��w��d��l�<����xaj���n����2��<���4X)�w��BJB.�kVv71�\�p�A�	b�Dt�w�WC���[K�%m�pG� �_]�oW�I2@H.u=�c4���"�@�3�DC�C8���`�a���2#�$�G�Ї��J]���Fn����ٹ��@X��P�@�P��� �3A���J!2�pD�\C~�`u� ]�L-	�=yPkPТOP1�	O���c���$�E�O��=H@$q�� �-ܣ4wm>�@����LB/����=[Dc�?��Iǰ�EA��W��X�
�T*G��ʴO�N"�F���fᗆ�V:�~�-'�Q>m��h����UÈ��C6R����?鴌�JH,���$���ø�;���Ҿ�o	��c�i�����M=�����|,��>c<���٧'��b���ؙp��-N݊�״��kF9)���M�"ə�(m�U=�(2a���d��	��.�<�3�cI*x�����^��"
�,�_�d��iU`CW��4��{P���s��� ~E ��� СA/MD�;Z���D�yy�k1 N�Z��f���0X��;��ҥ$��8�q�Vq=�R)���9jW2X}.�n�	h���/�;�����c�t<d��R�>Wj��C�B�Vy�S[��]!�j�g 2's��/�m��TCNRoI�K�PW[���G�o K�V�����Acr����g�Ga���6��&�����k����������Uz�l�8R� �9����C�t7&�t�5�Ɏ��xWdy�E��R�q0_��I��c�&�ʛ�I��
.QF.A���fL2��꜑>��]d���b�*8e����4:P�$$�=�9B�/Q��%�oÇ��&����@�M�F�K
��,�E�Q�S5�q�>h��B]�le��mv����AGHD\�e]�!�=�Ia�M%�(Bmy�^gHM��5h�HW����V��^�b�L)o�;K�8�E��a����AW��"�(��QQ����p���2t�=�s���%�e���g� �Q��<>{Q��W�Q�Ā�U�|��ֶx��Avv�� ��	�0��}��G��FBGWhl�>Fȧ���;���=��J}&g�?��&�Ǟ#鈾��k�Z��<nƳ�����]�	�,� ��=�:�v�e����YgX�V/?ܾ:|��m:�D �j��*�Yh��u�Q�&��KZZ����8�0�g"ǭc!Hdnt/�CW�.����7��7ɫ�	e� FZ�����r�!�&��ݬ�a�ԁKCݎ����c�!
�"!�9��t��3y?��T�y���]@
�+Ng�>�u��ziLɁ*��4>J�%z@�5MP��w-e��Qa�q���-��~�t{j_x{=����?�;u����}�2z0�䤳[��;��!����%�_���~���<n��-��!֌D�/'%7-����N��i�Oml����>�����d���f[{l���%/`���,A�(J�c��Y��jT����?_I�!jИ�w��T�������@"#0�T�����w7�"]�8c����]8,�E�z)t�c_��F���օ����$�����X !��wV&��K6d���C�T�Q[{�=E���P�T��~9!�HN��@�TT��u;�.)�K�2�m�t*%�aoN��Pk��:8��R7�I/>�G:1����C�.1k2�c95��jƿ������'oQ�+��Kd�@����H��NH��ߔ�>Y�.��b$�D��PY��t�K,���s��^`lZ�Yqy�K����@94�|y:^���q��۵��O3��r�e:{@Ҋ���/�����iZn@�yg6�y-�/B re��\�4b�|��װp���v#�!�_�x�X60��{�\d�|����fq@G���*sʁI���=C:j�P%�F3��iۚqrT9"�UC��0�^d�-I�Д��.�.���ǀ�ߟ���9oDQ�S����b�g�Ϧ6�^���D��^�:���x��8[�����zZ
y�3s�!ێlS����!R������?o�r{#��^^ڿ[@N�� 	Zs�4T�՞�
��c�n3?>Tg]��`W�A�ĪäB(��^"���pē卲��A3�F��R�uN�l�W�Z�	�q���/�vqRX/��6����*;��[��hS�-3�5IN\:�/�0k���g��� ��Sr��;��u4F���q�?Q��;-:INLN�>�8��iX}L�{� 1����:���A䘓��[��ᚿ�z�҇s�ŰHqSfq*���tֵX���G�/iP]���5dDD';�p�^��]���ҦK�Z�R����_	;�@���ꗡ��x��t߶`�9A?��c�S�&,� J8.�W19?�c9���'����V�'dy���{�.s#��{�|�y�oiYG�������Im 
{�J�Bd��c��7���M�@�"���%눯���[ys�˰�Zi��pS��oh�Q��۪YV���P艥*�&3����_!�PC0�k'oE� ��Η�6�	�@S���>����U�szwY�P�8w8�^�ʾ�ns�BVYW�ݒS?Ȼ�@�]�c6?���`5 0���GmT��+(��@D�6�y^�GUUaL�%Y@>}��.c�3�Ԧ�Ȝ#���r�O�WF��j�"-�/�!C&�Ŏ��\Wb�[��gp2��1�t�Q[&ȫ9�p%�n��yN��'�6�
���Q��QƬ*5�����h��U��@t���]>�>���f�����)�t2]���e����P�~T`�$=������!��0�#D#��nv�$���U���bjB�Z��F���If7��I�	��D4kX�o"P�	��w�T	Դ�$D���*���p�n�9E����[�ѿ<�'}y�!��y���\F���r3oʹ�����w��ʁ�Ô��XCGؓz��$1��dY�R��$f7�? 9Ͼ�ﾬ�Μ�qH�o������ݖ�<��i�=�%9	kqF�@���x�JG��t8���8+���g���o�JT�X^�+�<\sl��?'��y�DEd�n|!ۚ�^�gWF�S\��6r<
\8S>d��L�GΈ��)̶��L� ��
�#��&?<��߇TN&��U�Uu��؀)\Y�e��)/�Nda�P ���N��W����|P��^�e�
:�G!hח���u����:Ǽ�B���`B��"r˪c?I��<P9��r������T���X��W�>���'�k�p�6)��5�
�>��Y+$����g��g�Ԡ}0O1��7z�=�>{�\���/'����s�D��Hב�S�&�^�v��gWz�aU̴3>y !%�ZB��] h���}z8՟��gX�S���k����bYݹ\Pr{7z
���-�A�F��&�c]v��l��n�h�" d�4�ِ���(*-�%��|a�<J�����~{�tw���J���c})�����s��D
�q�����ܒs���0̈Z��g�c�>2i��r�渼��8�E%5�5�J9��8�r9c��QQʮ(N6�G2�dwJ&�[��l�k9\�W
dLT��W����g��aŪΨr��{�z;��m׮��?�"�] Ҽ8�_�Dh���s�~r�.+ޓ��re��cc�@U�6����ܿvҺ	>�1/������mx�f]��ou'�\5@bSvV����wQm��^v��nB�4��.c"4�[����m_жH�L������
��>�/Ά����P�0��^�y�{v��@0�t�0�Q�<��r[o1a{I�/�����*^k) �R`k��s�����r�.��;�r�b��P��S�xw�y��ѱ�-o����akw�J��-L�L@6 a�M?���U;;��9q��hcaG/n���c�ϵ-ͨ]6+<���?��;����E4�