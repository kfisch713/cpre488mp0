XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����b��]���[%���>Z�� �5��#zl�{��|�{�V�E��+	-�ߐ����4)�I\=d���z_UWN޸#�Zuf3� Q?v\7����xj��y���ǂ��z�w���,���鹁�rs#��WvVs&O͐��&i� �E�ȩ²U�cꚄ1�����K�j��d���`*���2�,5��*��q9g�v���1��k�O�lF�G�	jG1��"A$`컦pdK�Q�����,g�.�p�=4�X;D��ʗ����xJ~h�Jn2@���|��5���<�r����)��$�����f�)��qJ���&���5&$���)�7���FP� �@x������p[~ܦ$���2�m3��9��W�����a����"��/�?���K�I'���5Nj@po_2:�f�z��dM��I�Q�j���M��j���IQ�ƍ}��G�A21HĜyB�fT��~w�|�
�e����l�x�i��# �}	2�w����ŇnF_���;<Ñ�����}ŭ�!#�����!�9k6��+���b@�Mz�����1N�F(�؄	���ˊ��~f~��*s@��wD�T(����Ml����;z����w�(=E4=[��'N������W���ǿ�/���qn�=I�bɜX�;H0);������sZ�
���*hG]!�.�������+���,I�&�(,�	}e��W�|�2*ᡢ�W��	�_s���2
��>Vs=D��XlxVHYEB    3b09     f80�y������Ȩ������8�������b3��_=5�r�Ȁ\~�S�3�)������c+!���g�^|hS���K����%�RKbz��?�d�Q�bтǊ���5(�@%�H9Ȑ�&��L�\Lm�Ͼ��gq�t�?2�,�f�8g�wDc�O��ց��k��:H%�d{�n#�3W;�}�~�����my���,�h#gF�Y|ʩ�C�v�O�50pQ�P����d��An�[�>�tF,H6.��B�[� =���n�D�צ=��z�du��?���\�r3N�2�)d��j�1��<@�3C�\�b	���aE��d�'�H�N�oEAv�6zY`��*8B�?'Kp�}[�k���������j�Ӳ���!z��5b��3��z���M H0e�MI8]v����!��MuE����R�yL�Y���D���8�!�^����W�D-�n��Z����{f�2���[����~�f	{W^�^�	-�hR97��.�޿�W�R����jt�ME �����l{�����<��M�~��l�G�m�rs� 	X�5�9��P:�@}�j�T]|�.81w��*����?��/�K Q������	"�C�ʍ=�,c���a"�5v�ϧk�����x�2c��8���.%�o�����= ��3�:�2���ڲ-�S=��	ϧ�=�`�TX
/(XekTE��@�����M�9s�MȿX�|�v4F�&��\�U�5��E�g
Z ��7���+Z5��F��%�SY`q����[Bc�TFjI�%\�f^+R�-���B�ƍ���t����^+�v:w�Q��HFZoH����sQ�<�$��e�E�h3�|cRMm{C�]|S�K_j�k�h��pO�RYt�	�T��7@��+��\��cN�5�ՙ��0�bé>:���KH�I������ko�h�H�Q��;��7��$�;�<�y;	�`v��4l%	'8�E�_6���X�a����^�gƚ�ď��x7�I��;,
b�l��+]N�
:`�K;���.�#;y�~�L(6*�5?-�;�H���aOÐľ�7j�z��k���)�R�+'�Ĉ��LW�ҫ�n�]؎,����ϪaI0W��N�	ůx ���/=�i8ؠJ@d�GK�7p�y�R,� 3߬p�U����D����u��$Wu3����}d�%C`5a���«�e�մPz`���=8Qe�U D�+.-̜[�Qച��I,8+�[\ś�C�Gi@ ���nڏ�̛#O�b��2� ô������Ը�4\�����+��{�i� B����L��K�u˂�#�!��4�����0��!-"��(��Ww*i�cH۽O �<Qo��c�W�Ү ���i՚�ׯ�c��`<���n�?�ߖf�O�|vN�E��.}�n�k���D`�l��c����q`��̀�s,bKsL`	�xՈ��v�Ɋ��i9DM�OK��tȯ�u�% ���k�	3ܱj���Fأe����G���� nЮ��i����Ak%-'^���{��6\�U����=�U����$�n��/�/xYͺ��k!A��Ǘ��H�;z�"��;� �T���(�먴�Fj�Ø�&i#p'��U5Q�[3�6S*�Oش� a��f�Z�����3�l0Jv��g�hyr(.(Ǆ�g���}b���*`ۍ*��Vf��8m���ǟkaS��)C��Q�ÿ��?��:��� Fs�� �N4���_/I���S�\צ4�*[:h��,E�QD���F��ћC�.?����!�AZLU	 
�uued�V�N�p���)icHq�'�E)L�/o͑8Ȱ-
�����N���Z����5��]Y!M=�Vд��?�}d�e���lp�\@W��ܭ��U��M�o\�o�Oq�t��fM��"E��;,$F�
 ���)��j����Xt�Eô4&!�t��/���)�a�ݭݍ�\��W��Ѡ��q�#�s��ǺJtD��Xf����w�@�N=�g�1X�m��}��O� W���he��Y���\���;i��ߚ�Iuh��j���yԳ��tRJ�j���g��k�50�}�&{��0qޠ-����(������>,��c����5[Py6��Zpy�7�4�Z �yk�g�(�M3�����[
�g�������9���4^�3�=��.���l�f������Pn�Z��O�5D+=�u���1^S�3�u�+�[��<XB����	�?n/c���+$���٥�6�mLs|R�@�e�s��~R,�
�D�Rh�o�4��L��9��$����r�M��Q�%S3���%�3M�]�a0�Zۂ�3��v�c:�c�`M�w��7���<q-�@����Xk��Иl�6�o���͏�x�ͭ\is�e�" }��&>��%l�Y��Mt뜢��i0���ܼDL�5f\��qHI���cL��l�}\�#'�ѾgX�
�=Ozp֊b��P�*���s1�0r�%@�OVё�L1R.��ݡٹ˽��n[��E���z���r��h�Mā��kYm�&O�l�#�.-hAy��xw��',�%h�x)\V1U�i�.D"��T�BUpm��|@G����Z���t��()<W��L�ՈR;��c\iN��i�H��oN~�1J�����R,�8|Z��6�n���d�K��	q���t���ͧ��Ft��]M>В����k}��K��ź��ȫE�J�^ �����>�5EnâS��u��>n�wm!�ztgҴ����>��/q�np��`�����X-��z�3�_��Y��$�Z&�)�A-nw`�)�J����Sˡ �����e�\Z\C�|��C?/~�˝zue������<��g�Bn��֋�CƢ�UW<l�h.�؈J1�Pm68����YYF��jŃ�b	Ő��-��|-��we!\��T�	�1Vx,�ʦ�"k*��Zū�<�Q��ȍ��(q*�p$�+����┊������ �VCnk"�>�nƃʎ����h�J�3��S��?XeG�+���F{�N�d5�?��<k��S�D��ׅ�ŏ;�/�I6:{Ni��]R���;q/g)�*:u"׮Oc�:�&�,�36�5G$��G6�E�9���q�ӛ�x*���u�B���7L���l�G�.��I���6��0@�c`��u��r�5��	#HsL63�_��#}�+D�팜�CI��z�o��E�M�������:��)�ǔ���n��D�(��$̎�a9~���xD;�d���]���`H���\�[=\�k�"4q�>��f�'���Yb��K}�@H������-�-�#���%"�=<k�GoJ�]�G���^N�nv�دB���J�M�"�q�L�%e�������������:�m8�i��h$�1�e�atr#[r�x��$y�K��x��z�.Cv@7]�m����d��v�9;��Z��Y{�ɒK4��_jc�3�&��	?`�W9�N,��j�b��vB l�= �̢��K��E�S&��S�i�hP˪�FkK�[�c�뇯�`YS������18,r�/�h�=�M�|�s����S\���PnĞ� ��1�E�E��,�席C�@X}��:�
R>E���_��������i� f�6�tI����;^Z��u�����bh��4l LJ�#�ͨ,֣� �s�n��/�7��9�L�|"��;"8�`f;�.�pkt��x��ns�9�%9ZX���`���Q�@�qLl#w�Fx�ܱ��_t��Y������\�J_g���P�>�i����9s���U_Q�)�q<��o�����̉�#�&����C:���RpW%�2��l����n~Z