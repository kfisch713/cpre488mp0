XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��KyYR���P2�!����wP|g��r� qvq�43��{)����r��4\()�2(Lbx��嫪-�wy=F쪛dnV����T;�`������ꅟ�sd�,����rx�����Ɍi_Y�$V|'�z@�J* �Y�%��w_�=#�u
�Ȋ�`�2�L�5{��xǫ�A�M7~�D�?+��w����*��&up�A�jd
^����GNGVufd�(���#z���K{�g���sj�d����t6�3�,7�/�R;��J���lF֦l�t�F� j�`�3��A��X�u`�v��x4CDm�3����i|p�����bw��:���*Xצ�vX�b�{D FB���|���R �J�`�\��;����	���8���cE��G^�)�J��ø/� E���� ��'��ȆN�2�E�0"�#{}�u�H��|���w6����48�%�b�iJ�	�̴tن�
�&A=?�]�V��{��s��x�o M�"�b�A�L N�kU�2���u�l{� /�W�J���N�>k��D��Q��n��6�Z{�h -fs��9�~�$akig��*��1�1�(�����p�qlC��ѡ�������T��#0}��(CXх������pJ��`}�[��d�m�3������>�CmH��� h �U&dɒU���p��
 �&�<Z�k���v�C�C��~��{v��ս׫���2�5Pd��~��������Xŝ0��w��(�5`盷�ƛXlxVHYEB    1853     810�J�=�M�qً�����n��~�`�G䨝3�Mz})z�l`GЪ-��=���Ĝ��ڽ�p�h#ټcN�=�K}T�����[�OU������1!�2�%��`��j�����C����bw��)��@J��٤��⣷��:�*�<�� ]��uFǡn�����E.]uu`ǐv5zT
A�+!U�i.�0���*����Q�������l��g�.'�si��O���B�C��gG<�ne>[f���bc�\BYM�;ua��(���dp������`�A{�S3�8�a �3`1Ӊ��H�:|�����K̿Qcտ��_f��tCH%E��ۭ&H�N�3����v;}��ǫ�r��T��7���s�H3ͫ@�"�W�����Ꮒ�;��³���T�ܴM F%M��@�_�+�&�i��>�-�����0�	E�TG�˼�$��N�������l�A4jB^�,�_F����O�$�a���� _�m�!��g��W�<�#Y�
��3F�L�!�êU'�?>��T��~oc�*�"�dԡ����%)�y�Y���=H9����9D�f�$��\�}7��֓Sx��3"w��A�_�i��F�nq���;#�Ġ)b�Gkv�m�gڗ����)_חTŞ]<#b.:����!��|ncߝ�5�oNEJ��U�	�,�}IHR&����6�^�, ���#=H�n!���_Vb�I�T_�5w{m
�dal(��J�6���>+V�����0�q?�~�t�|��H��.�	ݗ���`΢V���!�Y����t�ᢍ�qS'�zg5�����כ�_)꛽��o�첋~À-�0*�`���zU��*������GÂ� ��GG0.��2R��
�P�v+4�?�.O� :��I*�U�W��7��G@��"̯T�h��1@"�.22(����ഺ5�l)DP�H��^�7([��R�6U>��s�)�OsՕ�5O�	�Rу\�iն�r����Na�#!,��k�_	}𑱥���|wW�w&�����<YŅ�d��
RF7�vt.�}�U�2��%����EO2F��;�CW�oʇk�5��{&�s�%���q��c�|�6*�s��lP�H��Տ��uA��a��Q� ��U��y��q�;ڱ�Ϲ���ƛ�C�K��i�O_����?(��%v*aPe������R^�	ٴ�Gp�=�L���$�a�$�;�I��Vi�0ߙ�<���`{'o'5,�/������!:Ꜽ'D�paq�%[�BT�8ݥ���&�I�m��PL�3d�����i����Q��K|�Ȑؙ=#��e#�� ӻL����~¡�|}E\_m m��7xck֝Gܼ�Z�k�
,���D\Иt�Ͽ�2N"�}|��u��1IcV5��9Z���j�9�Ip�
S�I !�r͗�E������(H��c\Ge����b�
���#�FB���Gƽ��@ђ�R��A��z����[_�Ȃ�C��)~Kty���%��drt��K��o��[�,�05�;�P2�3��I	�W����]X7a��,z �)�M�����y���Mi�E��׳./ؼ����I��1W���}�YGD�DA���$R�i ����ʽ��4��I���ǹ�=l��Y�atg�
��4�0�̓s4=��
�S�գzɾf"�+HSXI*
��w���#Y�|�Hx��<��~�h�O��BT� �X�ۺ�Fh7��y��QO��YL�d �o�Yj�fE��-�!ݱ���i���n�L�@jd�#���;Z���C�F���@����W�����J��[N6u���	��/��Y8�mP<SS�������~�v6<|���9m�;v��>�2�:P�S{���<��R�f����(�A�����l!���!�(�����#�e�a���^�m:r��'|g��nPC�0�d�$�W�=�0z����_����M��G^1���ܟL1�l�ۋu���+zIV~�� ��<(���H�-\��T��$ ! T���KN�a8