XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����]<���jN�j�s:ÉMl^�"�)s i���ck+���j��q�%�WɳpJ^�Գ`Ը�I\�#�5��X�C(�PhM���߽�߿Udp�令+���B��Ȏhʸ �u]�A��D�Gex�{��G�ޔD���ξ����w�������]��%������0�c�[q���'XW��)8"_�P^�>�y�*mO��}��pn�g�Ҍ���ci���Bv��D\[,���'8�t%3���0���/�Ҡ.wS_�:R/��a��a����O-���'r2)o[���R�W;��P���&mG=�� "�TM��*�r��j�d�\u>�32G�����#�k|1s+�'�b��mЕ:̴�[5u�(
�A�:hX��d��PU_�K�uޠ�v�xD�<pGl0r����d��q���G�X^m���PMu�w8֯�\�-(^�?d7$Y�����|,��5���;׿�"��n�PB��%�&qP���Oi�C��144���Z�Ȥ�$�</���<<q���4�QUv���^�U�*��5�4x��3���'7�>�j]�r՞#k͚ƾ�$��Њ�e9��pϘ]~lt��fʢ�BȖ�h�O��u2;���3��h,�b��|'>�o��L�Z0�t�6�5@�NF4�nm�q����s3�k���R���_��f��8�ϟ'��|��G�:G�8X�hB�2���
Y Uυ���ߗ���
K�R�j���Hzk⺚>��rQ���Ñ6ҵ��1�XlxVHYEB    3fdc    1160u!�	iT��#�?r)�13M5Mh+,��qf�CCDT�BY'�Lѝjt`\��$�1��N���'����r�2EAID9�w���Z{J�27Nb�M�D�����]��=��f����T�(~ك�fmR����7VD���ư�ja�ER7&���W۽�izB�`{Cĥ�c+^�:{�oD?DW�[q�!��N���W�L⊮��E ��D�d��0~m<*���>[K�p�/��OI-*3����l��|b�����x��2d���������-�j!O_A̠���kkt�����0�`���-��#�y[/Oaòp�I�\ٛ�1��7b�	�%�b�0�g�sm"�qK܆׀D*�=j����F�z���}	�{���Oֿ�.��5��.azr{�Tq�K�v
H��\��7�FB ����C���r�")� �M�'6��/�;�}%��������O�Cn8� �>�l������/�|e1К $����uC�'��-�9"�!�\�Cj�2��}�)76*tޒxt�l� �p7t'���h�0e��慝\��GU��~�"DE�h�Mv��G���-N���8��_�Ek��4'.MAq �^J��y�<WM�e5l��k�N�t_H�Xqy&��9ϭ*U�ޱհ�x��h�2is8�#�?R�P	R�aZ������=����.pv����/F����d(�3�T��1Ta��4�F�@�N���1�Ѐ��������R�h6�I��$wە7z���*CY1}�k'G���Đg�s`�0mm�������4Z��N7�9�������(�I�X-\�
����0muM�X�U̼Dl�����m�����#"�'����Eq����xyŌj�^hk����!�!0.3c����vT��(�:��4ye\7��I��6Y6��B�_��)�4�9��u���M�%���ne�^�2�L�b�y�#�1t᣻�U�Hg�[��z
��( k�Ļ��s ��-�m�C����.�cźx|�Wcغ���
n�pDU�����A.�6���Z��y(I��U2Klج�Nrc�w�������l�������	�˖Xt�v\��N�P@�����x�E�U�)����KWUD�Ǖ���Ҳ�8@Mh|���sp��>�;�+Trq�~wZG�o��`��.P��E2�����&�߬A@��Q�Y(^$�X�!C��G�Lˠ��@�f	Y׀��:���j��Dw.�����7�f�`
�N���e�D{0��:Z3+����r��.X��%�k�.���t&[S7��p��_�A��uL�V�ݛ~r�5;aPlafe�X�g ��=�#n �� u[�~�%����v>�Qe�]0��)�(��m��+QШ���bْw��%���~��Qv���^��$���;	e���7�z����/_ Zӗ!�\��vi!��k��E���;i�S(?6)�!!�B��^�C�N�������;�,΂��c�.TX�h�N:�qJ��"=��Q.Z�c/q��ҷsH޹BxYyy|}�1>�v�4<-V�����I��j��N◑U�YH����������mO}_1K$W��y8/篗?s�ǶT��.N��1g=W[�gkBPIZ^l��q� �;�JJ�}K��InC~URu���nvh��yOF�1��g�yޤ3c�~�2��t��HǮ�� I*	��B�6��J�˸6P�=e�)�ŝ�}@1��YNd���F�����￮�հ�ר̓�&VJ�P�����L��x�k�X�ş�
��A�A��H��k���,�N{։�O�	R�����\>Ч%���'d�D�S���J0ޛ(�58�W8���&gO�A)�քi�Q�Eb�uQ�kd�%���������q�FN�ҥ:�]D�?��g��D&-_���5�
O�JFP�#�N�2̔X�/4gC���	�` ��yO�$���I+�N�I_.�7�s��ɚ���{yّmF״5d�l&gy�l][��8x��lYݾ/7��KK�ϝR|F	��D�:��1鏂�dFr��7��u��@t������#�XY& ay��:6�a$������f�i�l�9�M}Y�W����
5\Z\�ؒ��2Û�T���I@�~�7��:H{��a�
�#0@�u�T18���r��i4v�"g��2�<掱{�J.=?���;�Ǭ��x3^����� ���^f����f<��Qh����[ۮ�PRj��.�J2lT�����߱��n/}�?*ﳉ��#���E�����B��"���u�6;��!��z�x�vz��\u�	�I����E�ܲ[���S>S�i�^3/�7q���؍����v����iT��7R%N>�6/W�u�"/J |TP�?S�W�J�7�p
O�qB�4s�\�d@xN,2>y�~&ը�&�����dJP�`~�Mޢ��7�����R���[�N��yT���j2'����h�<�4 �Աh'6%X�
�����@��4볇<k��$#�*ۅ�Oӄ�,�G\u��C�,d�#. (�@a5s]
x�y�A�܎Q$c���'���K�r΀�W�o�e��%f��K��U�|�$C�:�c.�[��j�~,(����ZWd�cp.�}I�Gd|i'��bSTZ��t�u(@N��v�q�'��Y1��9�̩�äm�Tv"�.���¹���
��&��1,��zxG���c��9���M`Վm
G����r�ط=HR:z�r���kK:��(
�:���#�X�aկ7�@5���=Wi��tG���O��=��X:ESA���Vy=�d�r,�D�iL�*���Z/Ȧ
�{�{��`��T��ƙ��'F�>{K%!��@�:�zǰ�+����CZ��&����r�OE���I,<,��s�"��rY�a�#^;a�T����9P��V�a��	7������b���5�n2=�y��<��+��Yi'�^,7������6l�0��;>D��_{o��(zN`2�7�W0x�;��-#g.Ys��Ҵ��,��'��P�qxe�}�o� �;��|�1�����=�aN�</�{y����`��H�l�������mS0c����깐u�Gy�鉙��Ƹ������W79 ~���ZA��^FFzT�m���m�{��W��� ˸��{�W�+3��Bs�Q۰ƺX>'rb�2�$��J�c�-9�s�'�F�7E��ޡ��=��3)��A/eK�n;�:��;��$}�4�_��6Q�$���~.p��o�+0�1��AEjTJ�1�)���[��H cz��0�.���KVXvp�E�6a.e0�uP��/����۷<m��N�3��U� �[�#�O���������,��M��;�c>Ƣ�㔅h1I�kgxS�v҂��n$��T�-�za�1��3��^���s�t���[?�����ֱk��tk�x�!Z��g��b8��N;�3�D�q�]t��j�U���9D\�X΃K��<w=��j�q�,q{��*�h���I��ժ;B�zZ<n���3=��g��
�����ߒ&m�%����CP����u����1����S�q�+7M����BM2�f#�F��dړ�D�K��?�1|V���ј�Arf�6�+�'���F��9��TP�]GɛsJ�4߲t	��^���$"����2W��a��=)�0��Q^�KE��Y(U��$x҉�-��SH��F�5���0����
�/.J�r��e*^RqC;K���N1C�U���/j$�n�7�r��7f��8�É��`�S,�I�o3�5̌#��Z�Α*�)�ӬB%[�
�t���@��ґ��~��G�6$���1���#�hO�g���>҃�\�3��H�FNb�|�R"5�-+GR��& �硍��UU��T7�t�b���~�s�F
����*�����?#�V��Y2�T�I��G��1���z�t�\a��YT� RN�{�&E&g�c����`��KY\2����Q����86Ai����!<D�n��l��W:��MOX����W��ؤ�՚3.�Ԧuoǲ�%�T��$����ý~t���ּ��Un�Ud�3?�/�NL6;�S���}ۣ]�����1N���Tmɴ�le*�#b�}�>}��7���Q��A�d��`;��N��3/�� /��^I�A0O�g5��)f�r��Q�qg���qI?Y�ǃv�7�;�����O0�^]'�*���L�YдD�ag3���)1t��w�:z��+EW�FqM�pF�:�g8�h.�č]�?���"w��S��m�M��ˇꬉ���@f&��� ���1�p���hM���bB�F�"}�ů���6�ܯUw��£'薊���K�@A���UQ�s�R�l��