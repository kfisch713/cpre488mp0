XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���reǦU�Q���u��.�ހE��Js�v�1?N�@c��b&߰�TX�w	�QW�G�X"�,�%���.�~Y�`��)�Q`���Ҁg�g��l4�^ʜUσ̚��,���&f��
N��-�[�}�q��"1*-��D!�i0�.,�� ϛ�6G�̋��\��,q\@�t�G��;�j�;v���p%�H�X��Խ�wt�,��0*D����:�9��Y�#�6��s[�>Dh�w?�_n����iV�U�aT~�C�93B y{��Z��ܡ8B�Y=L��c���v���>F�Gv8)�F�G��8��Ν |��5aI�_x@�!vJ��yx(y'~��Tt6�9�%�E'|���C��2��Y�f�}S����Q��,E��yʁҊW&3�X�4k���`�6b���!�U�S��)"�[���]_̫�e����3l?@Q
��] ���!uUߩ�2J��(��	|O��[E�=ôc��QR6M�`(%辠!�);'���7T�E�fי[��!�}¤`�Gg�w*�3�QT�l��S�~a�r��B�+� v=-AR���d�48���*-S�)r�i6�8�����$��x���*	_�T��q{M�sF�(��sb��|��r5X��N2;Mk�
��e����jW�DΨP0 ��4>�&���[�j�898�L'�ǥ�[��v�)]mϩ#�h�%@T�)H�ި���:^�R��ϼ�=�ِ��ҫ�㦓S���}�ٟNx�V���->�6���ꍓ���:�ܡ_XlxVHYEB    3fdc    1160���7�ʺ�m��Ѣ��7+�{d,ו�����������(�S�L,s�B��d�h[m�w��?k�O�-�$�pj�e'�k�p%�M�@���6Qj�����in)s�~�^�}����ƫ��_�.d�֚p�y>>m�,&�CN=�]��-m�&N������ז�Sy����?��)��D�8P���T������4Vw�ca	4�ʓ:����gs�nJ�2=O֎kM�ր�| R��x�T.���E:�}�Zx��fbwUC\�w�!ٺD�y� ] ���u"�X �k&J���~p�Cb~���u|�\n��'ח��SB@X������f'PE3�1X
H2�>�h�E�i�^���5KD�O�oI��W��_f#G��FjI���{߷�4 H X3�r�=�A�+��ܷr���?�'y �!	�)Ț��D?bZ�j[�Q2+���Y���{z濰Q���P�b:m�����e:����C�SO:f�	��]{�}ġd�BL/��~��P�ȯ�����_/�������*aS�@��s�����hr��jƘ��L��À��{JP'�ӡ �ủ����:��hE����_u������-H�̀�w�qѷþUq��Jϑ�g4���bۏ�o.Z⒣��u`tJ�����ԁ?[��j��da ���R��|(T�ƛuy�]��=tєD8�u=�B��r-�JY���/�|��b�F�(�-��k�t��J�b���d��sAB�$�&oYP�x�9UF�"e����JKw,�4��s�L`�M��]e��X��F4O؁�g�9�\D������\�s]؍����;+Ǥ�K����zm��џ�YRf�@�3֕͏��5�bs�0Aq�Y_K�1I�â�Wc��L������>l�V��|��-]��R�d����@�"�h<���"\7��>G�sf��=��N�嶨�(�u�@���$����Ȃ#g�KFrmCa�$)�	:B�$&!ϭ �[(�%��
Ɩ���ЙE>�2�Kw/��ٷ�rS�'!���<"�(�ip,�L�I�$?+Qe6��������>��-�.�-�e�E����6ݘ�X�*�* e�+�F�`�r	���>��0n�ln�C�o���[�@D�֌8L�����ZZMSYY����4��$e�E|�4-	��|�VJ�A"�N������f�"�KJc`j�o
�tn��g�'k�p��{K<�l8T8O����0�e��h���7�S�bV�_w$`��R�ʈ��'�dey9�Lm�B�����q��}�??{��t���{�v�m�R�<,c�\:#'��(�{�eqkm�ȈO2����WgC$�y�|�tw3oY���%�_tT^�v?�-����+)3P�G�I�#�́�9
 ��U@d����>R�ۯ�N�Œ���~k	G�L��r&�	�b�Cd�ןoYeRÊ���@�1��.��ӌp�.�e����_י���C�5в�ó9������(��|Tْ��р!R��C�gl���c�ݬ'K�/��8�b~S�q����Do�v#ƾS��ۭ�#-���}P��U��C�G�7X:�3���h�/�ɯ5��-�$�ؾ-�am���R-�KS$� ��x[�t�i�+�`�i����F!���7}/\Kl��ßo ��{ۍ� �>��zwF)a	�e����z&3=���F �:"n@uZ�k�~��Hx�t5D������9�8�|�xQN-ۣ�S��I�0(f��W�|:&L]zW,ZiYR¥Zz�vP�	�4 9�=[�/绍^O/��s�GBh�]7�����.D}']���e|�/O�:8�aJ���XO6���F_vϊޠ���'0��ɇUK�z])��eB����%_d�Ե�}��1����tٕ���R���41���7��-��/M��Իh��������\Y�y����Ƌ6�W5i-�(�%x��`F����cf��� ����;Q^�>t��7�,߯8�'��;�K9�șU.]&����,�LS�w�:��<[�h�f��9B�����n��7����L2��]�%"J��߸�(jV�^���Obg�ٳ��ȸ�1�!������嗲kw���1�P���lk����:���"C���,~ۧ�q^�2��'�}rX���q(�d�ž��Z���@�Dc/���:�G�7uG��*�C��Ǡ�2<V���x�D��# ���b�Q�X���glj�@>�;5�JH�
�՗��<���?�|{�N�J�#�f�ؗt��3��Oʖ�bct�V�s=����&h>���{�l/����K_��+�b�����
V��k���⭺�0a�ě<.O"�.Ӫ�;R8��n�Z��1�t9~�(�GF�V�sU�Dҹc���}����uzнYcR���Gl�����a�	@;��,���Q���Vet+2�?�Q��L9i6(������#�S!�������1]<ג�.�ʇbZ�j$�J�@�:��0"�m����9��{j��<S���	�U��cl/@^���֍
Ӎ�f	J��2��X�3��nd(�$i�JwY"���[ A�ȦK���Eh�ؿ\0K�b����f�P8E��ܸ;1~���FR�w����q�`�
@,�#�ٔ�)4�_8��?�Ļ���}2���qɚz���c9����mʋWL���~�y��#I#2"Q^�1^+15��ư���~�ϠkVⲳÁD�k�n����kr�ȭ�/pԀKP��t�$��#�ԅs�?�i�߂:�X��-E��E�b�ĉ���m(b�.�3D�*�T:Mk��a�L^�Y#��)��F�p�1
/)�����La����T4�=�4Ü��hv��=U-.l����[�i6U��.�������Vl�(�9�ZujĒT`�ǀ^�ozjX~��T���*auƱ�D<"����:����Y�3��9q�8a��Wt�nI� �|�M�io���n�u���4�fa^4ys�����Շ�������=Q�t������Fz�A�r0�pAd�28b�-T�E���H#����Z��2ˡ7Ye�N*���n�!�f�7e��&� ��ZI�`�_5ɲ�p��춥&K Y�h�i��L����^h��H���୩��Q0����3�3��7��d��^�Zhv�Z5v��f»=Z.�4i�!x!Qk��h Y���㴑���N��œ�����Tc�nn��edZn��%%걈Jf���*��Z��ͣE�W\�9|)�̌^RlW�r���EA��R��6�3������i�B��EM�#4h�7�ݡI�gւ�w��W�ιY"a/�Ŷt��޲O֟锆s~3�9��˶F��t�Ԧ����V����3&~�@9�#eb|'5�v�b�Jײ�
*��Qe��ҵg��{qg�&��s�o������`<��GEy1����Y��U{Ԯ��m��ߕ�}IZ�v��=��!A
�K�PT7w�*77�{��Fٙ���+��c<sc;�����=��ڈ����<��-�{�9�`vl�	�&^u86x)p��ě4P�g�X&鴚Q�ϖN^� u�0o ��:@��QUt�Q��)���L~��zCX���;Rg��v�0�G�dj�~��C�/��f��jT���֔�����oy�/���'���E���S}����*Ȑ#z�6L8����v���y�\�����,Q��@����0[���$�������Q��i����P�v�Y��)�	�G����'�r�>I��^fw�8C
Ba��T��@k5��=5x���B�ǉ�<��s�~:$4O��mU���{ڼGw�Pܩ���S���pc}��I��}J��J�PyoEr��iݾ�YO*����~y��'���9��ʈ�*	�=!?��ן�ke����rV�Z,�n-e���,�GW9�5R:�u6��/]�����H��G��F�O@s�`2o�!�����l ��٥MK+����A���K&X��e������~t�D�P��q���~�s7f
��lL��*��*���?�V�2�P.������86u��	`���8� �R���x�nY�hw-cl�K
�Lɤ֙ @�98�L��y~�g���~w ����(t
��DC��ְ�7�s������r�d�#ysB�	ϵa1zA�A�PU�_[��*5��U7ٸnv��M�Tۅ�ڶyeS��-.^}k��:sZ&(Q<W�Æ�D�*6�i}H��o��aҒ����3�Q���'&6%�Uu���Y}.�e�*�e�{�%H'p�R~�����	���1aM��(�A�5�}�V��3w2��+�<| ϗ�2�̨N��qY@��s����@��eu0uOwn���/Q�i�aؔ�����i��
��l! 