XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Kt; ����Q�K��K��^�ťv�)nQ)�@R�kk �H��[Eڭ��i-0I7�;��);,c)m�F}���@V��;�D<,��W'���wC�CG
��?���ڋ*���i�,���X]����N���gujm�[8�L�ݭ>�mz6��
~-|��]yk��p� �O^~i
�؉*u#�ϫ1��i�j�Cۓ0�-��)�M?�Ƚ�[���@�=�D�ʦ�#����c�٢��^6��(���M��$�5�,T9T�昇�2�@���v����2�D�ɮ�X����r�R�O�{��*��~� �	���{߂����_�,���W;��#11�H���u�@?�
��q�۾�=Z�·"��6{ۃ�$
��0%�,�MzY'N�c70�Ж��-�55�ټ;���ֳ��	�,�'|g'�(�o�����g����0��oԥ0��B�s3����0��P�?�`��zZwZY��!��/n}ךB�h@���"g��A��\}��:G횈�+�;0�'�+=!Ǔ�����3'�
r]�d�sF�}�����K�k;O!�@�;O\ �/�}� p�N��)�h���!M�㞗��CZ�gza��*�5�-\{a�jl���0���ZMI�A��HLXsD@����<?�� @�O�YE�B�|��@6䱿#+��0��4�)&!��j��a�����u�V�/�� B����`���o��e/���6�q���,�Q�T�it{���&���?|�I#WZ��m�X����}wXlxVHYEB     f6d     6f0	N˖�v�Y��G�7^B��5�b��۠gK��K��X�e�w0�k�a�?37X�'R��,Г�ߟ�K������ћ�w�'Ʋ�����x�m�E�e�JX�@���'7���!ρai�R� ��l��`dY��c��$���.���;�V�![g�:�Ǌ9v��,5&d��U#3�����-�}^n��"��0vr.�t/cJmI�V�!R@cE�	);��C���]���W����]�W��rf!L����ď���,C�Y�����%�3bC���+^��+\F���D�����PW��>T>�k��L䶹��X�d����u�r�^�^	x(L�`X<��H��9�JN�V�w��I׏��Ҫ���[�
��WE]��Ӿ���r#󌴢pEmw���v��k]�_=I��]I8�J �n&�J�'?,�� U}y�{C��``$<3Yz:`x����� ʸW�=.��44%��ڻgibl��ه���I�}^�@�Z�ߓk�q��U�t�~z"O����h�B$L���`Õa�F�)�&�>cX1���")P��om���a�� �ɦޓQ�nN�^��� g�%ɐu=������H��F�ҹ`M��h9
��;�ت0S_ـtq��&��l�6�!��W�UE�M)���>��?4���Z,<.W%�	1ʂ5�e�lu"����w1�����0:q���-�>���`��	��YA5�P��'&I~��Gc�[�Tm��^�P��%�����o��d��1b*+A֠�Cm�ul"���v+��>��
 ��Mͮ�%iX9��!���W��**)ڔ�&W��F� �$`�͏������E޴�{̹l��+�a��Bۙ�rJ��<��cT������=X}?���Z�2���;<�Z�o�lw����`���3 �󟉃�2�c�M�����Xy�b�.&H��Y �:��N1
Ji��I�S�½�/�]�)�fc�擰jq�F�ȴ��*QPs�uBN�~�v["��/�tvl���<����ʘ4b=q���c��0�x��f �����^�&ޓ���@�j�7����|Uz]Z����<�Z��( �&]�@C�? ��k��	��F��>���3@-���!6_���~��d]��٪ R��n�AB��2��D���R�6�(�{�+�` ��F"E�r�[��K�}��p���8<�Q�9$/Fa1�T��Gl��)�j������~ꠀ�$ް��"D��l ܿ��=י�שӊ$�[?�f8 x��\\>i�>\���F���%���N+�ݲ�"�E�	`��E;��=z�2F@��k�/����#��^B!�4�{���By���!}�g�G��Ya�O��n�K;)���B�Ih��A��P �ɓ`:N���>��N�����P���*Y2+�=��&�A�i��` ��1� �'�H��-��S�L&��&D��j5	�2L/of]l������V��g���\s�x	=.������~z�r��jws�tLN�)~�i�G�rbBĳ�֨�� �-�y1*{���w�kaRx(�?|� ���?(l�]gܿ���*79�vM�֚1�����	ҷ��`V^O4zytD:�U��9zRYj��k's���aa9�F���⩽8X�׋΄��R��RC�m� 4	�R���Mr}3��ї����w�n��gM���|�_*�(��T�}�좯�6�t��H�v���)�����oZ_Po!�Z��
N�;.�g_����