XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Z�E] `h�t{J��@�Bvmؔ��ߋ��?�^M��<0V�#qYw�3�_��׉�d�N���� �eNه3N����}L��pa�gqkI�\߉��`<)�ep���-�7���C���dL;D����n t�$�����v%ȭ{
�c�ފ.c��͵��1����n��pXO��Ty5�=Ol�F��"b��C�Pah$�����٫���N\�91@�d��D�"I>KX�g��sU�$��(|��pD��H�=s�,� |}kX[�:&>���������r�y[%m"	9�����қpj,O�tZ�ԩ*�$R�C�)
�k]����Vsz?��"~�K�,��5�bm�71������|	�h�畮'H�L&e�׀�!�l�%0]�S��/�yR�G+�U��Qmeo�"�|�i[�d�3͌�}s�T8n��}�{%3�^���/!�"��[>I�����Or�9B���MtW*�����F�c D�p�\b/�\)�AT�Y�����̭�qW�m������?�KT#&7_���6�Ub�
)N�=���K�ʶI������3��AwVՁ�$�U����J�����#׫���m�����>C�������ˁ;R��������;J�q����J2������{h֟��*^��M�OF~L���Mh4��|���L?���[��7��
D]�gρ��?ڇ�P:�*�Q��í�� 73�"�#�`��kWm��\IXlxVHYEB    6014    1840��h�`��4/EQ�`��c���I���@��A�9-hĔ�R�	n��t�i�F{o���F���ة@���&��0>�V�_!eJ=��J��`
_�5�0�.�畬S+t>�DYW�j:g�ƿ%/��p�_�hl
ņ�cHC`�?�s�	Ĵ��C8~�s����A3�͗���G$��0I����$�0�R�������h�,�Zι}ĝf��^Cg�ZC�����٭DK�j^S�TA����ۊ���z�:Ve�4��l�ky��ba�����-���J���Qq�WUUQq�?����#0�[��Eo>a�j��/F#������s��$Pgv{�3��e�f��*�Y�  �x�^ @�\a�v�[�rG4pinR@q�wk��A9�@�H��
������P����>eǖ�T�K[���0��F�u@��G������Z�ĻIH�*��p˲��"(�nd�9�$x��G.+�3!���c��v�&{|j�	TC����u�����;}�Z]��V#HaPUE2[�n�=�+��TC|C=��l�iհxq��ᦺq���E��> �Y&�(8Ni���V;�Ж��0�$��;S�"�73g�ͷ��ş3�������r�~L�����F�*���&��l̺P�He���|%R�&�\%��?X�RCP�8� �X���?��ܨ+�ѽ�V:[�@�O�?��e)pwv��z4L�$1��ǕO���jI�����o��[�!�EY�6J�c����1�J�R��A�>˙'�r��LKhi�Mnʄ,S($���X6�QN�X5}�?`8����NP��V����_H�d��������LL1�w�������a�� ^K������.S��g�����n=�g��о�:�6Pӳ#�|�����&�o2�׿�H�J�pǟ�$sZ]k8�V��µ֘jm�WL��5b��<=�ԻnSq=\�W BNw?�~�C	ծ�aD��N���\�x!���;�7���3����_.vxjfCZX�W4ca���lZ�ם�]�n�jH�|�f(���e6ݙh�O���]��c�p~�"�DV�y�t��9P���!V:�zW�W5m�gE�几`@t񬵎�Ǘ��.6F�b�9�f ������������fʴ��β��#$��t�-���,W��%�7����S�<��Ԃ��j@ƕZ�mT�ߡ,>[�b�@?E��$��K���E�.�C��++����ۻ:�agn�PF._.#�[6/'x���.w�>��j�woj:�������=��r�#)'�>���x���g�@��?b�*y�{+��7������ �Z�. ��Š<��W�>�̈́�b�|C�J�Kb�A����2� 3��=�{{�FO�{�4�b�¤����Z]�o��U��_H�Ǜ5�r���Ͻ���ܬ@���\s�BD���%/�*܆V�~PA!����9C��{����\C�Ibab.�LlJzD��.���-�:rS΋�H�U��ت�ѡ���}X�/6��ꍚAL�+�s!�����B&���v&��,9Z�ө)����?�����'1���������G�e���I��s)�fJ{42tt���hJ5S%8rI��@ʿ��<\�&3�����m7�27��?�<���J�c��X�|��o��}N�G��4E����:{&�~���2�1
Ј�#z��]|s2�Ш�=GnJg�f�����톋�b��w�e�;MUR=@�1�/���'<,�D�E9���b=4`��'�N?8��Ns�<�r������l�z�ZRX��l������?����愠�02K���)iQ6�d��P��B"eI"V�g�����Y�jī�ޥ�צ-��9z_����@Ӌ�������;��c'oZI��;��pӱJb>���f��Vؖ���1�)|�P��.K�HB��7���']ǂ�Tι����n�"q9�(�bG��~��ω��_R(5�=�(���])zI\7p4��L;�#jr֐�;���$�
Z�֬	��)&%ة�cV�='�����Q8������T ��ѫ{h�P�[�F�;���e#C(���ݟ��G*�y�P@Jq߆�U}��@��a;�͓p�Rhد�r\
F��7N43���f�&8u��7��;��A�Ӿ��rqG��:����h�>9�Ab�T��׳	�������χUl�gV�g�iQ�ziTg9�P��S�����&"�98Q_���}�ԑ	?j֍�u\���:�^�E��T��������╆p�8́E� |��A~��̈6�a6�v^������h�u7$M�?iV��+S�O��ʸ�B𿸱tF5�1��i\��e2��<�ȱJ�u�1�(	���R���-�}�:~�`�na���s��+ݩ:_T��'[Q쭚c;�v�8j�g�^���C~uvA�Au˨o����\�ޝ)����k���V�>�t�I��RY]]� �(M�Nv8C��6����]\Z)��B�C�c&�*y��z(u��D1"Xm��8���(�XzI	�Z�^!�H�!M.A\!�HS���숰#IL��ʅ�s�=k+�ڷ�a�T
��hn}1Y5���FGWK����<��^��햻�i=v�ò5ُ ��D\�G��j}6Q�f约y®�s$�Cr;�r]a]�M�ɀ�&)�?CB�0���",��'��R,F�D0Rv%5n���{ ������$ G�i�}���s�^H��Ɗ0������jX�a�P(������u߅$Цɶ�Я������V_��E�m�+��_�����*�����e\��r�\�$薶�����t�8���2��F
�w .ߥ�6�����c1Z��W|*��8%CW�N�o�D���NS5�bK�?��A�^���c�QŽ�_�vL�4 H�ׇ�W
�|]��	;�[���۽�: �3${�|"נ�rf6�4���~ǲ��J
r*;�j��&S87G�n�{���ɵb�K�;RC3��~�>��f&i�Y�N� 1�c�^�>���ėΪ\����iQ��|�ȶf&D�n	�>�T��nj�
xĭQe�]tx�����#DH�BT���R�u]��+1ꃉՙ_�|I|�n-b��| �����+k'��Bռ;�+���;օȳ���0��o����a����e�D�&�0+]3f��+�jsK�a}ㅦW.�u���ۚ[z���O����ܞn��0��R��{��� Q
u~�A,قbXJ��l��	��$^2�h��G��P#���ė�6�}�s��P����I$+�`S��OF<��"|�@H?��
.H��>����W��۔�l�E����q&��G�/��\P�o���j�`�z����c(��2�<���q���g�p)\�-d�]��{����@O��?=���[�!9Ӊ�໛��H!�*�F�TQVN��H L�/3u�!Ъǁ�,��QwiINo(��kgQژŒ(鼭��O��K6�`���A�Ud��H�R�ӎ��[��s���ܲ�ތؽ���E��t�a���WdRT��_ݦ����Sh�X�ƿJލ��qі ��+s�Uv�hZ;"ra77���������@��� ���7��[X�7��]���x*�^��u�k|�*,J�C(1$�V"�jZ���'�x
 ������0�~��`��C��ʤ�����d�Y�<�:Az>̇���`�yu��&gB��2A�TM0�,�!~nķ�]���Q6q�C1����3Oݞ(
)��	X�R� VR����D�Wӳ��Yf�ڸ85[`�e�"�`'�y�E�q%v��^���Y�?x��Ӝ�`v!������ө�ᄌJ�����<R�;���롙2C5{|U�1%�A��H�2?�g������a���7��T���'��ޑJ�R���f��^"��d�y߱�<���Kwv���tw�U]�Ֆ��^ι��� `ߜ~1�=��1q�8��[�]��\J5鑽ۼu�ڂQ��5��j��w͵�)CY)���HD�5�'Dt��7~2�4�T�){���3�!8�_��V�\(�h	��`�Dh���ψǡ���^���j�ץD9�I·cW�]�~N��F�5�+�_� &��ő_�1�� ���.���8��Ӿ��X��61�ܳ�$�x���	C"�Q�?Q��k%c��L�_ɬ���!���~��E-�Ewc�-���s�����R���9�T OS��ec;����v�#��GH�qNËL5�|���{�iz)S��
vآ�Py�(fD@D�rZ�-�_� lB%�X}<M�҇������bƫ�����Uό������I��� �F~3;9[IVp�i�������${ŷ*�Ӵ��r{�h����
D~S�x��(��g�i�2&�.�(K�
@���KeS�P�||*Ύ�x���� ��H~<ْ����&�+aJY4ۈ|cW솞a���wv���X��4z�^�Y�h�HW�bρ�����������w�h=DmE�(� �`��샿@���Ujt������5�3>R��3�M+K����-[�rׂ��;����9�O����h��e�4�q?e�K���bm�ڿ����Q��LG���@�.R+3h���W�8��
]�-�2�2r�ˁ��F���Ӗ�E��G����c��PD'��2.�p$�
���������R��k�.�i�#�>^��G�V��R�Ϯ�|��SI���C+p�)F��dkXk�8~��� ���z�_��2z�!a��m@�(�΄-�m���Cjʸ�B<Ë�����>"	-L��B��/��oI���7��֩�+Ƣ��o�N3rx��#�jw�bΚb�i���cۑ����m� 8D2� �$ �,d:b-րLDC'�~�E���͐ A'm�t�LC~z	\{y���Pm'Fܽ����5O3��
Tq�L[�B&����_�_����\'���ϊ���W��={�S�Ru����Xe0���y����rZp�.�"�(ٚ$�8�c,v���#ea7Tga�Ѩ��}xٞ9�Lߗ��~�L�����H�瓞��sR7PF��v2����߼^˄����8��ĎH
��{�/���u�_Ne��b���0����X��~sB6����m����+��~j�w9>�,DJ�e����xˮ]��,��Ps��7<�HX��~�v����P
��|�c�\��ؼ����*�(��+����s2���!�	����Zuء�]�����\)yȢŽ��]�\�d��;J�	�c����ޯN�Zf0�*��K+n�U�Z9W|aC=/"P�P�G���'�C�!�v��f��=c%Q��8pWa׶qC�]=ڛʏ�f�j �{XD�' tDcY��|�b�_FA��\�2׍�XE��ЦƖxdq���r��SS$��cM���%�p����B�~�����N) /���Ό�����
�f�(5�rXGy�A!цw�}��}�908k.Vֈg�AHw���`_���G=��37�������u���-$�_f)�;6���֓�d�}k�%.7�x�k�W�g|dj��T�k�c�3����7�)���i҅	S4�7,x(`Ng�4�u��+�v��f���	�L�U踨��*Ivf%E�,�pȮ� �^��Ck�
BH���1�*ϊ�i����ES�,�F!��a����j@�S}�ϧV�,�4ࣼ'm�IG�$V�O»��c��3�p]���=6# ��I[ Q4;���qх�pS[�	{�ï���z����H� �d|��J�(�zS�3��{�'�7"�,k �~P����i�^:c�5����-�g��F˧}R'�H@�jyw����s�Slc��#��Aj�G. �ɇ!4�1i��^���g/iG������'�fn�啕�@wK\v�ȭ�(������$���=~�x��/��e��:"�l����uEZ���؊����͌�yHh������!��y�Ujj��E��ރ��ú3�8b� ww���V��H�o�)$�gN�.��O�@�7�YU����h����I��#l�(CS�O+8s$*6