XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6^��r?��9-��6�_NK<�3�{�K��Q��F�W%��)|�-���7[�=�Z�4�w������|��O!V��$�Q;�4���㕥��fU�<�az�RҔ�S҄L��Ґ��o��-��(fqE��d��%F�%%�hքs��&lrpc�{d�tN������f!�ܝ}���q�9��P��WY�q̈́g�T����p��WK�:��1�(��c���2 c�F���7��S��*����
���9	���\r�2�K>��'��[�+9 㢳��E(���{�V>�A���k'����u�c��pHL��l�5׻n��cgG���	��XR�K �!��U�r�߄=s��Q <�[YR�09@3ږZ�C	����~�%K�m��L 3Qֺ`�'�&\�v������`?�Y�B�P��#�^%�~�ҋ̭X2�����|WXnF���8��p����h���/*�1�4���P�
E8�L��:���`�$�Ds�V����j�k��R:�z�I؅�Fzr�K����m�|^�XXD�9��݁��G�]g`���7�7&��ձW�0�>����I��*ds�����W���S�H!�s`�������-b�O�y��QU�b߬�R9��=MY��_��Dv(��Ai�P+�'�a0v�gvգ�*��h]&zW������9R���e�H�0�B�UWJ���T���f��َ~�&����o�������'?!�v�9'8�^!&��ZKXlxVHYEB    6346    1790}3�3�Ñ����E��r�c�v�eV<wò��ϣ��	T�G7��z�����)4W: �q�� ���0t2��NF��[�s����V��G��aE��`�k��2�4Ԛ1=��S>N'�߄#�|}�"p�\�Xa��&���
��]��G��Mb�dRW4EoI^��(�1P}���<�%F��R��39��sHM^�z\�g��l��_c�¸��%�L"�i�����Ҕ�
���<px�i�RðMw�C'�S}��Z6�i�T,�d_��{(zT�F/�5�F���Wf�6��%��wwl����<�H><w3�=Ǎ�*����_R�a���=� >� RN
�0�Wu/^& �C�ē9(�
��ϺE�@:/�Х�};W�����Y�Z�Q�f��Z#�?!��I,��ϓ*�V0>� x]�0ݩ&��=����n�yU0���&���������ۨ3�茶$7(�fژ����b�j�o^[4)��2�=����ÂQ�+SmM��#�X>�+\q!�hr��dהg���� �m�B�tv����"GMS�X�ʚ�,,kZ��0٢}���QK��ҟm��rM�K�p�"��r�dXF��ouq�J�$D�LrGaRq4� ��.�Q>���"�^�ă!��-�_]��p���ޔV�~ p�8�{ն\b��:�jF�?��ۆ���Sh��5MB��~Xx�dKQs�!��0x,�ϙ"@���qoԖ���9�)էi��J9�z�z>D�w��FCz��V�\N��vp��f��y����@C����A?���^��n)��>�O��"e,1�c��&	mԓ�:t�[d�C�*Lk�J_�o/y.�2�̷C��
#��*<��uQ�25.��x?��h��I�1��qE�L ��u��.~�nY��f�ݩ��+�Ӻ�6ߖ���=��f��Q�����z��x20���[H�ô=��{1��w@��o�tNQF���,:@���`���:#-'��9a��7��D����9
�h�É�ĩs�q�ea,�oo��*
��+��W�b��76o�;��̺�/#���&RӮ�`��thw	g���$����T�AMm�㖌m�}�8CJ�ͪ�Xm����zW�A����{������.��j8�m�.�=WI#6v2�|���Y��|8�IM���I63�TMT%�w��g.�U��_��\�ΑS�`���du~.�$�==A���y�x�5 ��ܿ��sX�~���`���bi3a#��L�=��ъjO4u���*Ô��d��,��Ze]���F��+��_�YE��
Lf%��7�?OEJ��S�D�X��j/E�Ti���2q�1��M�s~V��>k�!	-�������4к�
T��>t/�/G��z.�.<_��N&��	8>[6�� �*�Op�����=s\���4��5x�qw�U�S�V��2�\��2f�H�[�44�+�n?@|MҘkƯ�u�3������*����-�^��1�e�7����4��'���
�4:K�p<�=E�V���+�Kg��O·%�1��1�X��.]��`K���<�u�V���b墐�`�vL۝%�b_@}-/���it�wu�U^���ɤ5c8-53Ѐ��b�7����
�(T������a;@Hm�&1�#$.��ng9� �Sd��3�����26��)y�`X�l�2"o�<K1R���[5���w��>�3��G�{I�1�����+Z-��7۳6�U�Z��f�w+�-n�I�^OO��];�y+#X�=�G�*4%�^3H��X9���΋���-���;A?E�E��'����
�f���lѪ2Q�=zK5%q�r����>^�v�N|$n�Bf���bZg�Z�K�1VP��"M�Y#�J�Z��s!�C�xM
ɍ<�ն��Hi�Uc��P�5m�q�z7�dU� o*�A���r���m��H�d-d�y�胇x.�c�Y"��Dunh���(�;�
�	�Ի�2A� ]�G���J�E�Sܜ�N���v������5�xa��/� �Ξ ���e�9�
��H��ф�rֹ$���vB�U,'Ƃ�g���C�,�%�z���������8�agӠb�d(;�����&w�{[1Κ�!a�㵏g�' Ǡ�hQ̩]�*N��l .�x��z��Bhq^yL��I��-�5R�|���H���HA)���G�zK�ˤ�z�d�h�����ÔFo�k��}�QT��l'�� �z���`"^�����oWu��=�i�Qj2p!�e���>��[��t	~m�/�PE��f+���$�a1Ͷ'$[�<�h���4���xo���J82��!��)�Ҟ��!���.蕰XQ��2��G��(�M,e����Ei�z��������<�L��'S�+��� �٠'���@�dY�)0�أ��b�D�'�[�*�������_��g�md5U�̢u��Qg྇��lxq9'v%'Rm#�ڦ�-e����q�2�/MV9\��S����ܵn�?�K(�}G&��ҬLyl�7Ȳ�;�j�<ԋdF��Y�1<�4#k
�#�@��C�b��  �Av/[�yv.��2ɔe�2��f���ʎ|� c�����.6(C���ۊr�f��|���U;P5ғ�S�-*����Cl�|[�=l�m������@=}(h���ԩ�A��o�h���`�t�ʔmqc��A*���(��T1�u�0wp,&��t�5�8�D�����U�s\�5�W���.}+MM=�=2U[��)U��(��h}�7��sY�Ydw�F֞euxd+>�&в�?���橝�[	\eu}��Q'Z�z�ʏ	(Zr��� au�Ϛ����~��j�]l�F��.���+)n�KW%�kU����ec.��ެԕ���k�����·r����b�Kx�ΩN���3��]�Q!:J4]S�"A��~�d��(�n��������U{�EfEG������R]P��t�=r�����b[M&�Uw�VS��x�H�!����<i�-��P�7�����V1���Zq'��L���c(���4e,{{��l�3�?h�u�|V${�Q�R߾dAO��E��~f� ��)���BF@Eccy��<a㾼��T{��j�� �1�v6��<s��B�u����5T>��8Ӣ��6��:�3����_��3�C�����,q�쒱�s��t�@��;A�6�6U+�H �\/�9$�Tۣh�`�p���W�[&uh�L��E�g����4{a��l�ås_t���M�U���y !�t�ln-R�L�.*���J+,�yCZ�I�g�Ё##�p�￠�R��ʵ+�d<�;��)�{����-�7ٳ{+���f�UF��/ٞ����oMz)�:4{�:�
+�7L$1Z�n��WY#Մ�%�O�/��t.yX'~đ^��s�>�/�3�	�ؒv�괵���B�݀������p
�Y��+�냐ʷ�N��t�MR�[DeP1U�#���P
n�y.���v, Ұ^e��wt�\��*V+��4���KS�8e��g��A~Ҩ(��%�Ŕ 8��p�W�� �#k_,�`�*{�ϼrG�Ccb�kT�IZ�Жj�_�2噯�E��b��M@�)�i��mR���g��92Z_��Z�?�ڮm'H�������秀y��&�ɑ/3ll�P
�n�J/���4�������N��O�}�9B��H	�M�#���V'���P$����<�̾��f��Ai�x���go� �/��!�Lu*\{�(��5�ر��c� ���Y[���[�'޷���V�T� ٮqc�H݉�Yi�+�
��d��˓Mdk[Qˈ*�����T��Y�����>D3)���צ�-�����M��s1.õ7��y�,�GK�YX����A�<�Q�z���=e=�M~A���l�S1����JPE"S��I�}=�R�"#�(�n4���~�`��"����=8\SFЂ�:8e��@���Ђ�#�~��J�}�m�. ӌCr%&43/n0N�'�0Bkq����:wQ<�[�����;sWT��v\��d�9��}Yc�oh>�)��KTޏnoĪ�����·&5~�q�O�p��޽x��]�H�f���3K��%�p�<��R隨V.�t��.�T���,gX�/�����֝��4�@R�.fw�?�#�q�Iw���H�r�]�E�K��������;r�]�󡳵�ո�2��[�؄!����m���X~�c�b������ǐ�E��LF�]������ym�R&�;��D�!�z@��j�;z-�bd�!�+��GT9��$0�p�&篊�fKl�o��?�����W`G����S�'���*��j���4h �^ėcR,r�)Ŷ�}n�=b���4�1���F��'m�޲h��������,S�F��a�s��$273w�+�z�A	&���_Q�RƷ��e���-��:'�C�Ҩ$��x�]�mf.�sޫ���]J��1R��is]�.^�u�s~��H7o��kq��A��O����ttӷ5�I[:x���0u�"���ռM��1[%1�l9�{������py�?�kWX����@/������h��i�aJL�h��ߐ5�mR���1<�="ʭ��{0dU6���{ѣ0�T�۲;i^�2�q[�Zg-y�
���5����B��w��ͣ��FOWz�z��d��8���vG���G-w�������UXP*
�:��XH*�uj�|Z1���D���Q�"�l��L��S�g�fC�B��%��%�Z�
.��o��� 3��O�L����>dR���)�׀��:;8v;������0f���%����3�.E��B4��;�N�)E�Z��g�V�B�֥d�A��q��UH��'&%���jL<%O�d�$�,6�g��b]�"/G�q���?��<�^�p����v�i�������l&H�0U��Q�&�D��5����p�j�G��5S��7�8b_c���EW�LM?4f!��c�%Q�4ׁ�Yؙ	�J�˄eH)Hl���P��N�3��A��4�ќ�yHtڝ�ϡ����^a��IǛ�gp��C��b3�-N�VWC ��e%_V:c�;I����f��G�<+�W��uw�6��w����<�-�NR��ф���З
u����G���ML��k"���njA�<0j�н��q�;
�g���r��]�����?B��ցo{�M���w��¥fLdJ�R�9x�ס������%�:sCú|��I���|�6���Y��P��J��F���1'�1�}8v�E�N��Bg�JҨ�Fsq%�L�� ��_z!,ǔQ'���p �e��ތ�
'�KOo�|zg�'1_T˾<��km���2��}�_9�O#&f�!#�Ă�1ފ1x�&@�[�]�p���Mm|H�*�%ş஽��(Yu(=ؒ׈�xD6�ˇ�l>��o+pa ����GA>^CM�Pw,_?Z�Mu����T����BP;j1gb��Bh���VX^u���u��@$������yu_i�M뿩������z?Nl����tM�נ�f�A((w�VT*~�υ����O\A���9�u|�������'��M��,���h>|*���6���ܮU���x�9L�oǁ��i���r�7d=,��+�ZQ.Ί���<
��&� uX���ҏ�ՠ^���M�S|����yC�g�w�'͐�p�!��;&M"�Z����)\Ye]��?����k�aX��(��(�0 g�w�Ə+�8��ǧ����N��XH'<��#F��������Ї���Z�@s
p�ȟW��	(O{T�8�4�,�2�i$�����'�נ񡁴m��NxX"%@u���a���&q��dE�̢���@�j:c���Wf�s�`�;ܰ|�����X|P��G�w;�N�>�r�F'S�22���J\��'�?;SSR�h�