XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����X�4��:U��G�7��a?��.���8�%X�lac����x+|����s��` ��3n�1���+�v5���{���BX��F���J��NvEh�X��2��Ob�A�#�l�rv�� ����qso��'Sz:���	u�@�H��S���j����.�}����
UK�&���<��&�7��(@��	;=�	B�I�v�=E#I��Y��n�vlG%�L���i�/FR/OEN���R�_4��O�~Pಊ3v�7��Sl6��/����x�U}D%9$���}��Z,bU��t2�9�0 �[�Ae��[��hW�V�͎{�k1����8�&�z�J0��vE���1��)�����+.���eu<������hɞ��K6�� e�o���F'���}Xʚ�Gw�Q��H��7�Ԓ��� �;ڕ���~��
�:�(��lSԋ���B9�
��5=�?�wJ�ܕ���0`4�;w鑔5/��\�@������;�Ew:<l��~2���#�ɒr|�X>�I	�T.1>q�n���?V��(r�$�@|@��O�:��,�CMB5��p)�g�p`�	8�i���[3�}Ջ|;���{ƺ5nl/oI�E_f%��Q�ڦ��s�5t������'}��5`:��8Y�����KV���O!��5��VGC�� `�3~�&ư�<�']|B���kF���b�pz��!y�y�^�X�0=�8I�~�h�L���w�{�ڼ{XlxVHYEB    a037    1fe05Q�z$R������!��;CQ����}�^�.������eFզP�7��'���*&�/-L'A��v�+R�V���E�w�d���q&�c�!pq�W�2��!k�ذK:,����6��%;��x���.�$U���.�K�����\���k�.��Q=��s܅���o���طi!�KE!�FU�v�p��$Q]�tCc�����xV �_&������W�JHW�+sHLrβ&@&H���m��Kױ�~j��k���-��6}�������GRc,q��� TL��B|k�%@
�_(�&��yɭ���а�s&�he�ch� 7�5Fx�#A�m�62V��`���f����Iyɏ��^�c��Z��еƶm����B�Ys�3[&-����;�G��2SP�:�fK]+.��H�� Lɪ�5��rݡ�`���L�Ȁt�T���Z���l�1i�.6"��.�i�@K���ez4��L֨�жI =KW���>�j�p�iٖm�֩A������*e<z��YW��	���&���c�|4=��烊��0�����Κ�V.��PԠ�YOD�t��CQ��p1w>�,��I�!�o#̷�A�y(1}��Aс��a����7
�{�_�W`�<���He �{I�[�!��BͻbWhŔ���>\Yk��>f�E1U3��~2�M�=�$7m��հ� O/��֚a�;?��C\��/���9xJعb'�z��>Ae�V@�>����0U��_��f.����aHg�Ԑ*�	�:P��3��%�Z�Ť�K����NW���Hx&�7/CW��o����������Q�I�c�y�{t�[�BS�lB��}
�%>9���=�"���/:K|�C4���ψNB�E�ءs`�x��`�ߺ���6��]� �v�ǖ߸��[�'�:9�:^k�}@t3���r��.�Z  �%���r�	F�d�u�h��T��zvm��Q�@�v�����ӻ�&��tv���.���ml�&���J��G+�~��^���k"���P���oݎ�$e4z%��k���G6LU���6���G��}bx-ֳ�g:�ii
�]��Y,�����Ģ��^���]-��vIٯp�\?ؘ�P����T��ׂg��?�N_{T�����:���m��5O�]�
�~��V4_�� �m����D�h��$t��CĮ��o���[�(�z������n�n'ո����X��s���qb�B���L�䀖C��$̶D�/m��������P�� 4d�K9���_����d�-d$���#�B���$�	��w�ׁ�'����
h�1���S���
D6kl�S�%4��XUs���r�k>hę>`k�����W�ҍ��^E�V�9d�oGe����R"cW������sǀ\h#�%�Ӆ�l�������x�Lq�<����e�XW��)�π"�E��O�A/*���vK(�sJ7"����o#[[^\��m����zf]�rŕ ��?��Jk�ّ`j6T��q�_��w���:���mt`HV�^����vE^�� ;	�4��?�ð&T�N���2��t���A�,$��q�#֎ԗdcq���%=��U۽UC���D�؊c��$>����I�S����6��(���	,L��P#W���|�"ȗ�m	E��Y��CX��- ��K���>����^�Y�k���lL��l���n�,b�1�ܤe�x��W!�nA��|6���%�N&"|T�]�w����x�C8�!��������QZ?�q��<����.
�q���@<�2��ɯ�WrU}����P(?�^�Hu��}�(TS���n�j�,��P��1�kM:����Є�#�k]�U�((����}|��Lvb��5�}��(2�����yX�Jka��zZ"�w��5KFy����6>��9<�	�#Bp]��$���e�n�u����ITB�g�m��l��D�MhB�%[�z������4�?�(lY�� KpI���t��?�z��>u�@���&��Հ�Y8=r� �!Y�W&㱎��BtF��kG�{��k�v�	Ϸ����I_UX�E��n�u�ʑMifd?��AmX�*/�_.�r�����K� ���6���9�0oO�ث�Pc��P��6ۏ�{8�^<���� �_(����7��������6rX����:afY/�H��S��'{MZ|��-ԗ�ڣ
+~��l:�bIr/��}�<$MJLk>�o!3Ջ�_�E��.m9�L}3�R� �s���$�t������:=���u�0B�_5��k���X�T?���#xvb13��a����e��;g?o⮟���0F�v?���鐂m=���S	��A�A^~*�+����n��BG}���
	9닰l�N�c�G"Q�s�G2�U��zBpc�H���o��De�5[Od���4�f˯;����p-��\�߱;���cI���e��}I}�H�8�����U�
���)����L��W�أ<oR�B���@����X%.C�ͤ�*!�۫�����q�����;|%3$K∻��JOy#�)�ˀ������swª�Ffr0�<�� �.�2�I<)�R#R� �>)-�נ �W>s;4�����.���Z�T�T�-i����Od�}��tP}};�;����vp2�cL��`�,���$��%�G��>a����*��i�+�f[��������4(�h�Q��0�ZR	k:I��G���{UK�}��cM���-�x�pjEJMd���y�����4��;A�F�Y����9�������n�o�l��"��Zk�s	�=�s��T�Ef�ѱ"��ձm�K.����A��# >�Fx��#��I*����ܔ䖽�7�g�X���M	�ЪY�*�9���Z�X)�o9�t������.)]kˍ�P��-u��qeM�v��ޚ���lh�og	���b�V����Ħ:��|B��G��� �i��/���nIb� cKC�Im�?
�~k�f�(�d�2������[�\�zA	W$Q���Q��z��ؼ%kӦJ��&�i:��ww|}JՀ�)���h�͟v�������\��ī�����];Nkg�O	��P4a���Q��F�팆�����}�7�ǖ�6G�'����.� $m�$���9$��f�/
��Ȃ�B,�\cłc��b�i�������g՗F#v4�ʍ�~���4�s<8udp�/.'u ~�\�9�8���BǨ3ŽyL�T�^��|� Y�����ŹC
�͑G����һ��`1�u�q�����¢�Ҙ�.��x�y��ۼ�Ӷ�f��mg��'@y�c�:��Ug��Rjӵ�Fl��ګ�숭�ܜM@D6'��,����ZܲVL��#V�N>r�L����A^i@Dv��x���S1"��n�^�뉠�`�]�fk @�� ��Ɓ	{e��k��U�>`n�|3�.�X�pJd����Yp�W&��4X����6c$�h�[��L�؎�^��l�4��n�v�q2Y��Lc<��i~��5eI�<	 �riQ��J�SmWЃ���*���tJu$#w�9E�8����]n������FX"�H� A78�����Oc5�eN��[�GE3�v���)��}��[1(QOJ���j��Y��c�
��9��X�[0��e
�|�i��VP�.x
�3'��ك�����%w�ʳ������3�?�Wݤ���𽜃�X]'H�O��Yp��I�R��ICO>}銉/,>j��6��>�!;����td��L,�>,��3~mC�Rb�~y�z*/U�������M�%u[��Dsțh�X��x�Ƌ0�b�A�Н�_{�w+\��:�<�`���!H*C!�\��M�j��a&|Y�R��ݱ%�do�)*��d���L$ܙ�˳ٿ^�a��Ҏ�tO f !N��V]���(!PD\�&����&2{D�G� Lۀ�d��
�z���"���Dh�O�>��g�w�A�ԙ������;OQ��GdΌ�h�bD(%�#��{�oRN�����v��d4�v�.����r�V�f{�]���Eru�	�7q�$��[>V�$�Y̶�'\�Ý��:
p4 P�!��&{�`Z�f}x��TY�� S�څ�{�:C�#�H�2j
������_�t�t
{��$���3s{I;�[���}�al���ɣ��}eڒɩ�z�/+�m���Q�MV��F����c�;�mT�톼�<U�����&ݮ�,��!��Ϊ�G<킠}f�S?���+�9e��,��\^������w���.�ꩍ�,��[U(��U����&-�߆Gk�4-��KU.��������&��a�MǓY_�2�Y^�^%.HӒ�_d]p���eS�[XV�Q^�ñ;W��N`NOY�5D�vM���p��J�=B���9Vˣ������ư1�ā��p��_�x�N)�2ǜ�V���%"6K;œ��b˺ 0�h�ʠ��$7�m䩶6�g<auPݪ;w~�G렳��g'o��fȀK�Ӹ1A�w�Q�$QAM:��S���9=����z�F��K�;d4-�Y����� L5��(���ͦ��M=YG������K��fA^����:�-����q�G��W}��
��d����8��T�������:����̠
[���dJ����QP�8�a�E�w��g,�����lg����W�dk1-�S?!��9F~?y�Ѳ���H���#ėE��/b����&+V���(R|qo,�_пi��%tbP�.�C�cM@۾3-�!DR�Qԫ��\*G�N��^ǘ7F�{r� ϴ`y�x]+	����T�����ã��W8�b�����g��5>\Z�w���e� V�RQX�����CElt��ω		"5�4������"�Ζt@�Y����aNV�|!����[�~1OBf����<����zD���h&ʝ�9B�z��3�J���]f�m��I>/�2U�J������q)����&	_�af�W�AN3걓U�D���ץ���A�� �}B�gJ�ώ�*�����yN�c�%���[Pv�h ��T��'��A�oZVY�7�x�7�{O��$��	��n����]\�����No�ѽ*�X���k*̧���m�B@�qt$�T-�$�UZ���)�/=F��E:�d�MP�@	&�XP�� ֱ�V��k��A���?�y:�P����2��e5{ze�cl4��(ЗH};�m��s�|:&κH9�&�吁ѠI�m���^=������H�P2�8��i�%�L� �w-���#�D���H��U���LZ���o����bD�y�|��m�!�]��)wW�����|#�@��Y�~"0�s]�7�y�a�wc����o-l��&�ވ��d����}e�oa�]���O�w��b %n�}�D�<n}_b_�C����kW��SmB|H�?I��[_3�Ş^]s��9y<*�߫Om$V��<��W�e3�:➣Q���Ox8kp?�<v�<w�g
�+�rO�9�	eD�1c�L��j�W��h��
^��y������=���L����K�+ņG�&A� "��A/������fN�Y��YCB�2&~������`�� ���t:6�
�Y�6�<;��D���W��E��i�n�s��������>����U�b��ط�إ��"I�}�ߕf�VCڀG+s��jprH6X	�ߓUu�g*n ����D=���'�M0w�6-��+-J�>�H
�	=;���wܖ�p�ab��X�T?�ҷ r\6ۚ��P�������� m1����B�tr��jm"A���!�!Op��t,)ٞr��gxt��)HF�s����$/v2��_v�U7��s��Xŷ�P����&5ڃh7Ona�f�]k����Jq�4P�o�=�'k������]b�q^�+���<
t?��24|�E#5&s�V�x&O�Ǥe��g�P�"�Z�X��ʽ4e`'!Hq>.w�J�@;����=�t]���*3$��ߝJ�6c3z�(*<&�%�%֖�F]홣���T�H���6����"� ��>��K��c8��e�x�o���
ܷHi�����wV�䅃��a
��3�c1w�V,"�����s��,�tf-��h:�%���z�2$���eT7�aԚ�Q5��NԓӴ��;mYa�շ:_������Q��ܬ�WXE��9;�
����pX�m���𵲈���E��~�?�h�wo��d:���p
�_�,,ٚ������� B��d�4/��j���qv�1�S�ҫ�����&��Q��  �nj�����A���HE�C��] ���x��+�	�[���>"�ە� so�v�t*���ӻD��E��[�(�f>�N��U��2���F-=߈?�&αK��U��n���J9���D�,̖2p*�O���EI����4M�B�BU؆&�X4؏T�5�/�ֽ�â��-�����I;�vѥϽA�w�H�Iv�'W������W^L�Q�"�̟����f���ֻ�����FO��.V�v�Zl�>���HiRBGY��.~�bg�+�g��N�9��Q�R���!�#���+J&����(�M����	���,��[^�r/��Ӊ��Qޥ�nP��Ml+l�U�����$0bކ�ZNIb���� T[�?G��@N-�7��S�S��^l9����8#N�;��¡�]���+RS�+��C_���s��n�h��)��s�n�A�5q)���S���8�E��*�Ҍp۬a�gXC%���Bѓȥ߄^��r���U�1� �ƽDt�,�Fc[�,L|��A�e݊M�z?_�h>������R[��;�9��4�1��%n*:� ��0ǫ��kJI�)�Jlc�豗 k�$y���pD�ĺg�p?[�= ��[w�0r���*Ĭ�J/|У�ș=�Ni�	��!Rg� dQ� ���K2�i�/׷���"3"pM.�hJ��⸁/���v(4�8�l}�{�6��Ky�b/?;���L��Hui�D�Z��y�綻#�=��%s'�$�ݬ�q��\>�V@Kz���|�L1s��{��6S��w1�ʫ�{�^{%���]�7��c��V�Ў�p���Ȳ�:�H�6[H�P@��S�dV��/;!��D�=y�$&���CC!iU��YDwӮ%��AAP���G{kLtf�w���wyy�Z;I�������˔�֍bC�<��׺�^3Ȩ$w^�G���U����q��a�F7^X��ՔD	Sb�#�N�t�.�'�d>�\ �o�Q�����<���ԟ1� ���+}9���0��n?�n��sc� ��<�ڃ�����8|ڃ�_ɬ#V�d|0�%S*�MD�A��%�Q�%��ˈǛ�
�l(H��m���`&վ3`f|Vә&T�
�j�X�C�ڶ7W����A&����4JOomʽfɟ�Ub1R��6W"A ��`p��H�h���6�1�P3��gVR�����=��иJz�;[�W@ �EB���O�G ku��,�䁸/E���nSZv쿓<���\�(�s8S�p�yk�i~
L��$�:B2�5�۪i�R�x�W�?�h���+��#%}����pt�6�>�=�����N�6�C�ڰ�6�nv�L��n����Z'�[�p�ig��.:��:�'5U���H8����!��x�OE�����s���3%�.(Q���Cu�fJ���=����{��8���dw@	�J}��Tt���֋�O7$���0�[_ܸU]�tj��c&��|+���jr�	(ٓ���Y�d�L:�'�"�p){�E�M�����@7h3	�<�Oh�Y�	՚���gf~;�n+>���Z� �����[5.�%�AԦůIn���,��E(q )֦X+��)�l�P�,ݯ��@S���/����ǯ
[,vV蕥�m34C�/�ѵ=��x�