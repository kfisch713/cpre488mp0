XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����՟|���1����G��ip�p��h>�����J1^�(��?;�9��Ib�z4���UX�4��x`�4�(t�����y4�S�	���	�LP9����t4�� �����*�4S#d�匜HF��qxgݰ��7T&�h*򡍌t@o.����E
+�g��6<���R�^˫��T�%3�g!^��L���gG�$���9��"iw��)5+u|e3�a-޴�'��"�N��{{�_ ���oL�b���l.�KW���Ô]F��8qG{�Dx��z�u�D���)'�%|^�;NdCs��q��OB�U�$M����Ǭ�<f��(�vWx��3�;��{lf�phbg�x}�!�X`������Kwズ�߁
�u�WI��>�����;��&^n��?*)���B���^V	��ZNcU�Ƣ�p�iCBP�Rqs�ydC�J�5+����kL�e煤���(�Oٶ;z����0]��	��x>�C�c��CeBtZoL��$xވ� �E��&c$���=H?jʳ�D��r��oT��=.$�qګD\�|�2��F�i�SA�pu}(#'9>I��)p�<�@�T�������(!�^�����,�ėZ2;��˫^磕�pQe�0����ǥ �{��95/EĖ�l��̧�����d�.��a�K,��#->�(��E:o��t�I��������W�����q�If�	�L�ø�۵A����З� � ~�*��J3ۄ*,��.�������|E)x=H�3B6�XlxVHYEB    42ae    1110�Vꄡ@uL)�[��� _r`�-�]�⣵�t"���מ��Un��|ܰ�3���$Lu�,�����T�n��=ns:��m��{?RJ�X��̙v�����P�h����̃b[t�'��K��������	k�v�����1������L�z�Q�chj�i�.�"k��c뽁z�ѡ�d�%P'�f-�M���B,B�c��E�۸c�Ɩ��gp�ٙ�r( y��~`�*-�U�~�$������V�ݔ�)�E��B!���/Gs��;�����Q���@\�������j��wZ��Y�8z��L�Q�i�vQ Mr}�OIr� �n,d��DקpU�e:�u��V��h���O�����b(d	w@��7�M�GkT�>	�,�>���QK�?V���9㩣Ԕ�Dh�2
�}67�<@h3u�������Ӕ
^�N}?�sa�)A����Z��ZP���b�ؠRB� M�s��q*��t��R\Z�"4�5�tI$�bb��U�g��q>���q�����O���xgnM�����g9�Is��&^1��R�`��X�e��/r-��R~��"C�_W�,�)�4�9�����4���0Qɿ��kp�u�S!��]��>�:�;�x$�_�0�"|��i�lEϜ�}�R��avXS��4������E��WP�P �=���t k��p� �j0����i�*� ��4{�)_�9��j�9
z��p|�aT���f=f�P�Ԑe�75X���M"�/�s������ٷ�!Cj-�F��)Y�"_m�
Gr�{:�4#)?�J��M�(�o��h� �͑���g�z��6k�>R\�${�3yG0�.�=u���z������d�x�����ߊ$�j���*�\��a�OBY3�����J�^pe,���c���Wf�`���wƥ����[Iz��U.ڧ^�ۊ�$9�٠��j�v�9��2��	t��������]]��A���m.���De���\�cb��/v/
�oe$�)><ńQ�Z����v�>�#�y�1��ġ�W.�L*��U�v����q�1�=�����P����t�aq�Y?����R������ߚ�F�F%Z��o)Pc��v7�1�,�툗:�ϯ��~ipԉ������i���k�wx����T(����%M�@�-`3�

UgbƩ|<z����	�A�?���|�~�$K�<��雇d�,�ۢĴ���ܸL8��e��>)o����j܁�� e��:�����	��3)v�c*��k�� R�ߦ�ϣwSW�`<P�6Ez��:������G�4�}.L��=��Mǆ�\��9�g��"�6֡R����� u��3j�.9$Y��"�&�v5��W�Mш�aV�BA��}
�c����qn�.�B�焝���C|X̍�&p�\gM����@װ!��j� �T�R�3KQk��ȴ�oj�e�j��0Ū�T��4����#b��/S�_4#���Sf�m��/./v�E���@~?��@�V���b�j�ڋ�F������o(���",fv2�)�7�5��_��0�Ť��W�FvF�������T��/�����8k���x��W��;	S<��W~�/K0�H�o����|IfQ�T� �{�����gx�}�ů6s���B���[���X�H��j׬�T�ƎΨ��?#�\��q����Ӎb�9�, p���s!��.�_5��-�dDJ)�ȃ��^H3��CAAoE3B�>^6��;B��xx��f�K�7&{@s��zuB�W��������#��5��q��#Ю{_A��G�R��*��E �]�1����&�����KJq��C[b���7)���ȍ�u�ӆ�a6�R�<x2 �{��zjF'h��{��N\9��>�� Cx����
��� �z����嶝����7��ධ�����d��-��<�iO)�n*h���H#��&����2!ꬵ�n~��p͑95WDl����P��'��F9w�3�&#�H�T�PfQ�
��P��@�x�yɱ�1G�J���{�F��Z�?1}�"6�� ES��Ʒ�����E����y��;*?�����l6;ѓ&L���4�Ɯ����I��|�gV�7g�MӺ����h���'F!OK�E�j���W�����������MQ��p��w����P!����LW_��t�S�>��}�����+�沸�
~s28�D��f.j�6�d�+p�v�d�ț�3�s�/����h�XI�V�7�g�7��x� �U��S����E͐�7�d��H�c���C(���~�:em�p�yi3�rL=��
��3S?O��a�R����eo*Kf
d��i�$2����$:�K��Ȭ�� �E2��̜RȕL;�RG\׷K�?����ܶPe���L!IXEUdZ�A���ϫ����,���ћ�H�&�vZu�T�M��#x	o�i�k0�aPit�������-ep$�]�K��]Wi�����:.����V��KJ����٪�����M2�~*�V-�"�/�#h	<�ɜySV)$�]`������Dڜ��`n�>l�@�(��C�us奺��y]��OS�b���`#L�d<������0H�Q�kv���Bs1ّ\�����$7�vΊ0>uPep�t�)T����b�+4��|���lHÝ �l��wi�[0W����7�M�I/>0�°�\��:ܾ��{�R���p�}�Q.�`���z��wb>No�W�@����j�]f��剁��*���ϑހ������gK�5,�O�/����3�9�pa�	��m^���89(�9L����Z7>)���U�%G���|�1����$������ߑc��T`7�b���rbY�-;)��!�ױ���$��5e������qѹ,�����0fq�a�����k�J��T�̣�uϞEs�u��O���j:��'*���g��Fy�OX�Qar� �����r}0>H^=�X��O��.i�}��r>�k�����;=����%C?b�/�jGp�mj6�-v7�E@:��;�	�[�/ ]�Y�<J5�8�~��>�pYs��zyi^r02l��Ƞ�S�c��mUg�	E�t�u�Z�Gk��Ĵƻ4C���Z@�:K] ��R�JLge��i0���ך��ٽ��6��=�ú~�"�w���\O˘��cq�f�Ӱd�����ȟ[j���8
�d���,x�e �/�b�Пvd6�Ў��(��󜍑>c�w�F��i�1��'1�K��LM���7pԁգ�F��$�_]u���Q� �@=��=�|aL5�SN���s/���Y�:ubFN;_�<��j�S�SJ�����> �9gֻb&�Y��*�?�JP�^�4�1���b��Z��
R��
M�
c}�#�MX��F�]vT���0�R��(h��a��)�Z��1��Y�%�h�����4F<J����NĿ�����!a͆��GR}��gP��&�o�:7�1�2	%���\��^%)W�4�e���}@-��u�F�u�Q�s���Dө�Ά
���UX�d}{4�@ʠ�L���8��hgZ�1N��3g����YwJ ���lҔ�bV��h�W�B�M �fE��QE������}�Aѩ����٘��#sy��D���a=��d]weNCW��I������IԆbz�k����}�K�0�{����+�p��Q5�=r����^:��eTBg�YW�+m�5`���]j�c�t�8E�2�S�%0B4�����?L?����Ā/���WQB{�ٸx�e<D;/�j�Awn�l��Q6�5a-U�23��vYjh�<v#�B�\Q܁�bU�3��ȯ�ٌ)Ak:�]+@��R뤨���v^�t�X˯D��}�@0���62 ��R�w)Tτg)�A���>#)ac�l�B(o�L��c�nGn�K�t��Ө6�eh� �ia����h��� *#tTLSR�4�T��|Dt�X;��SR�FJY2dˮ�o9�',B;�i\nܚH��)j��ɧ�V�k[F���0�x/��Ia�%�*�' u*K�Ze42LŃ���æ>���0��4�r�0�	�*�L �e^.:���F�`�~�R����}C�п�ĉ�B]O��qw��1)�L��?���h�ό��*�Mw ��DN'tt3�|�f�����^��%r�֌�[� ^��k��QSD��n�qH�)�S
'���!C�{T��&"�i�]�Y[��$��k!	���Z�~<\>uX���c|>