XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���e�H��3�oC6v�w����'IY��9� �CI�s�1���DX��|O��{��f�]��y�W�����U�3�o�:�6�"�8f�ȣB��)�`��}� MP�8�2IVF��)lk�B28���t�n�A��U��Je	U	1̴9��
���!֋3�u� Y��!�ȷ}��7g'v�AT��K���|#*�4��!o�������P��Z ��Z�u��H\��f<�l�c��{��K�e��GH��:��F��tR�·�ֶ�ޒ��V�u$��������.�s�Dc������v�Z�,al������5�u���#N��'���V=L��'s;�<*��~�{�4V�-8�̑��[N��e��<�f�W��U?d/�(^�e���+�]Oztb<�a�� n_��M;�{{Ǻ�l�!��`��=�-�1IRm������=��{�g�B6����?VY�ͼXG��8�!��a��X����S5X
9W{��݀�~z/�+�n��(�o���KК�-Dқ�Q�g����c'�PW�s�9���@`���<���c@��&��t�ȍ?��nz>F�w���z/�X�:��K���L_(O����:�8{��(-�"�>x��ҷux�T�:�r���tx��5�1��8M���x� �f��Җ�"m���Bā��l~'����$�8qߛw?�/�y�;�`��xI,DzA3�#=��׉e����E��:[d��_F��s��v�s�2����ï�Ηgu~���XlxVHYEB    3b09     f80��A�i��v0C<"������g�uU�ޚ�����o�dQ�� ~)U��J�M͎Cv�]?"Je��V����<�H�G���@5|02��S)�X�3����D��>�/4�pL������uĐMi��'Y9�̐����>�z�!�_�����D_hF������S�9�u���}ۑ�4�w��9�B%Ut%8dg&\K덀s6��&Qx�`S�5����.E(�S�B1@I��׌��қ\c놜}p3g� cc���j���?~�@`����R�G����[E>�[���K�m�IvN��́/0�0�&jI�n��L+-�@���E}��G����}ˣ$��jb0�Io:/�c�!�|��H����������k9��"��qwO�I�&>�v�2�Z �R� �����W�y�$�..�6��)�x���R��
��=�X�-��KCe$�m��Q�	������sge�����C��j�l ̖vЂ�BX3�����|uj�$���@\qCH��)]�y��v���J�1�ڣ������S��{9ESm�GE�X��\��H���U4��׸Z�c��L�U,t��n �)������wy�s��`��>g���Ჽ��bJ���N��w��îB׵]ܝ�XQ���6����O�9��E��П�e���;���^Rk/��s75ɪG��:��6 �����@�U�r�pbAvb�y|j2��ɭ�Q�9�b�Ґ���S����8��3����0I��$f�S�=8�x�(%̅�;ArC3�'S��+�����qFD��{+Esr�G^	
]�j�;At�cz�g�9j)!�	d��o�8olrX���-�N�Nl��u~	"B�"�l>��7��3lHL7t-���е⬗�M�
iL�M����iFU[#�wy������Z}Ҹl�4a�=��?F;���=�����4�b;�����8:3�ia5%G���>�/c!�D~�)D\ T�i}�a�f` g�[2,�٘�|$A�|�V��1u �@�8����Ź>�ȫy�3-����mWDg��~WQ�^��o����m*+�	R����J���Z�D2��쏗����2R�ō�TD�Ay��b�zy&�dp&Hd�V�g,{�8v�J�,m�5����d!�"?��<g����b�L�@��/�X{^����s��ݒI&2���3���������l�ݳ<��mڨд �a���;�I��0�XB�|q���挈�8?	$�f�z5���~�-�}`�tP�����`�K��lY��`BY�~|"��ٳov�\ baX��R�Ű��J�{$m&o�����ԗMC��;1m4��l�Q����ޓ�B�>�L5�c���q�+�UWX�ޘ璟��tȆY�D|�B�s��5�A�2u��2@� T�	Y�q=l�T]��U�]���Fz�qg�h_���Q��b�f%�{�瓔#a���|�+�3!=9�l����w�K���NșV�a���p�Z�^�Ғ��8{vο��0�KR�Y.��)��=�=;o�u۝�cg����v���F/���^���q�r7XE����=�?��q��pCf�����HU)Q�2>I@R^��C�$�$/Wq��P]%�0���'8����\2,�@�=����Q�:�"a:y��I���n�Y�[1#�>��l� ڦ�М�*D�[�����O��<y~�\/ni�d�oay���w�m�V�X��缫�l՞���/3J�J�@�S�^G�ZU�ƹ���Oa�0_����w>�^jn�6W�J�kFo} �n� �������$&���]�����|���v���߿�����[�$����n�6�<��I���.�)nɲ��O��; �nm"	�Os�!;��6�j��R���SYO��e:]�)�����Jh1#"w��ַ�¡Z�����x�ٶ�vy+G�+p3�:趃��-�.��Iٓh�����U�1�j �}����>C��g��Ň�0��w�S�����2d�Kw�I�_tk�L`��zp;�>��},l\��X�a`���@'`���Jr�y���Nl�j�Ɗ��X�3���:Xw�@�Y�LN�U��W�0n��я}�?�j�@$B|��:G�?C������U�(�����Q���m��B�6�m�<36/�&�5?�l���wi3F/T�W� H�s�%��e��!l<j�迸����q8�L�|>�WA4m��1���v��+��;�����\s|���ۦ.k�C���yP*����A_ͱ��W��ZoNickMy׸���7���h|�i���=lU�v}Oz�m�zS̑��V1�{�m�<1�|�x�d�M��3	���c
�c^`�����v-|������	&�����v=8���٫�� ������X�R" Jˏм��*�Rw�2u��=�H>J����l؂!�A_ZU����~���a���L�@��=�6v���w*Pɗ���(�h���:B-��	Y�;Z���s�j��jԪ֖D��<_���i>-Z�f��I#����pb�S�SP��;=���K�_�>8ܭ��x��%B��NwU1��$�N��Z;�d�n��?� �E�Iw0!S�Db�E�
jIk��f�w�b²�8�FN�W�5��R�to�*k���zI=Qg�D��XA����'��Z�,�	�x��P!�� �pC�\�2��o���D^���ܦ}�;9�"�S�V��>L�>A%����*�(-;�͗�U.�'�~��tGS���9s�o7���hΟm1G����5uh;�d�$���ET�mW�BQ�"��T�X�r�a�*��i.�w�Z����a�(��^�v�e�;;��~����D�cK���,Y��u�ag�1������-�_���.ygwn�s�4�9/�P�{��qkgc{g!:1/�;t�*.0�+�lԏ��m���@�#������,#�����~�ve��?�:nn%��*��)k6��'\'䨎�.j� f�"��X)u�56^X����[�̐�Ě�|�7��KCk�.Go󮓽dP�m��P�̳C�&1)Q<�X~�W�!����ؽܺۈ�C;R��s�����O��e����.��s喠9N��Sف�~�Ybd�����S��<��I�{2�N�`����	b�Dp
AX__�'0��JIGB�wߤ�ظ��3�BX'%�J5明-T�$]S��hE;�Q�3'��:�S�X-��f.��#.&	x"V�綏7(�]m�t��`�~~x:�y�$��:X���}��{�>vXyV��5��.��X���$�
%:;�����pg���L�6H�a[�?�(AWL
���}C�Ÿ}Nʇ7���G�pMd��/8�k����ht��[@�َRR����x2��4�.gļ�����<�
��	�*o�R�&N4ɋ��q����x����~ٍ���ui�V�)Jx��S��d�?$ �W�{ۃ����O.L(���ܻ��=�M驅���K���	,VJOR�**��՚DU�M��G��Çn��ܯ��=���`���·�3ڠ�~<k�@��PS��B�Q)�v����� ǂ�EInR����_��e�aS4M��e<���D��*��y������#M\&6�-6Wr���K��%R��N��^�Zđ���-�	_i����. 9����h3�'��Ҙ��K����'�=��/ڿ���Fd.��]�U���a������_�i�``���!�i������9X���!>�8+������jX\W�Q1WΘ�O�OZ���#.�f���2��3Mi���������P�j��&��G�r!��>	@7�W���>��5�fͫذl��N�+��t���>b���{�T/��T�_ͪ�S1[/�V1X