XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����F�� ����""Ѭ?W����7�,,��}j�ۋ�9��ys*H>D���.��j�84�R��ͨ/ƙ�_ut_��N$�l�¾8	S���ƭm� ��g�G��=���莌�Y>��	���{ �U��%+]�X��k�@A]�'p��@�E ̤�Tk���������%X=-�2����d�J�Yro�C.�t	Mi���z��B�A�j�M�E\D�\+��g�'�ѭ���ڍdI�X�� �5���t�o�=z�M5'�@�f<㧛����C0���:i[a���g�M;��ݵ�r��;�.����
/T��3��кL�[ﳶrGD�g��bV����׋���\}fJ(��p����ȝ�Ct�^
�SVP�˜�*���?�,Lc�����Z|�q��P� �ڝ� iDǯ��\���\�x�z��V R4f?���,h	�T�Ą�T�PX�R�i�����P�ɭ}��X��L)��h�u/㳪F4Ts,O��p�\�Ř�Ma\����1+�=,@"�}l6fO�2�Ka������5��ń���R�7ϲ�i�ŗ�ꡨ��zBh�w�6�{�l��<\�]��۟��E��O�`�rC�f���v
���d����vz�r��w򍡹�Ĵ�������s�b��/}-pm��h4��M!z��%K+[Nnߖh�2�+u�2+����O󷱃IU���atx����)��rz� aݩF]�8�4lգ+æk {Z�2F�r�esXlxVHYEB    42ae    1110���7��^�q"x�P��(>����,}M������o_�
�cDP _~Q�L�]� 4���!mi��$� o�6�fE;kZ#�P+p��_����&���"v�U\�ՇřE�!�+��������VB:&峗����W���M��îy��K�H����������ѷ����JW�
z�ȬVBD\�F|?BiZ*HY�u}��P|ʋZd�Ko��?e�kcE $�x4�W�������̇V���H �O�w�~M*+2Bc׸�* �)�II�y�@�]IՒ�P���Hl��Ñ�aC�aǬ�9��G����Wŋ����ן*q��0�����\UF����1!����|o�hH_:z�������ie�k� sP����!�/ձ3�p`��M�Ŭ��i���G12L2ps�OZ߻���n��o�è|(�Q'��:�2�Ԩ��}5�kއ]�x�z��Xt�o����}Rs�š
9��GQ|��Xe�� 	I��Ш��Y�ճ���w�E�3��%��J���_�ID��F�yk���M��-1n�Kz#3΢d��E��g��{��5U���r�&���^�2�´���̗o�5R��DX�Ű�Aj"�	�P�\�����Wۉ�� }�b���K0�Z�O�U�ɟ����L�w�yC�P\$�<��+#�['��1ha���}��x����A�莬��]4+������J���Y� �M��$�n�%3�k�[+�mA�#�1�}��/�I���V���r�-ƂD�v8�
3c?����]��z ��N���1�k3�Ȟ��Sg��LM`^�q!��?r�\���.�%J��Bu�!W�n�0%=�y1ȴ�X�����.� �����:��V�!i��.� ł��(Jo}�z�n���x��B�F�;iA�LJu�+�( ��s����7�|L*�耖L���1ܤ�l@UV=�%W9c6�����1ˊ]uv/ddx�j�j���@�NB����-�N����#}e^�֑�T������]� ��q_)�u@��eX(�1F�^^�*���WY�܏�ٺ���ߓ2+���������sG?���Ғw3�j>�&h�=[�Mb��1��婂N�h�k�	4R*��oLJ_\��jϲ����^1��V�*���T�9J���]3'����5!IQ���E�_S����O���w/ U����d��/<*�)\�C�
����$o����H�!���iԹI�`�~h��>��?=]X)
!Jj�� �!<�2��`&D~^�뚘`o��у�B2.�ih~š����mwao�$�T@���9�5�Zuy��F��kl �y�gYD�H��,� ���!i���%	�H�x�,!g?wk��v��a�3�~:���3h�� V�_P��r�<����n�F���Vz�*�!��Z��|�RN�B� ���\Z���"&�0^��[	+xhSH��:�>����DD��0���!��G�fEsM�_? �ӏ��^9������/l��O]�����!W-Sv�bWy���ϓ7�jll��ڢRf���j��E�rX�g8�HF�a殒��NZ8����^������"Fء*��.�w�����2�W�}�]n�/(��DV�P�54,�pY,�L'"U�#�F���k��`�=��}��@�R��$~ꊬ��lPyh�#IǢ�w�O�G������
�`!���ZV)�s���x���(9� sF�H���׊
�f'����G)P
`�1�K�FO�L0�Lv"&�)�|E'K�E~�o����#�@k�Mq`��R1X�!\��י�¤|�ۘ9��+VGXe���qﯖ�'����)�/�	�ۛ8E	z�bsrĤ];�b� �l�̃��J~x�˃��e���.g�O(N͙d�-W b�ZL1�+݃ľ�2%�Ž9����J�E(0�])�����-��3-.#�U�t�|����]�͚���� �ўG�QmE�@��Mf(���/���[��2W wzA�	f`��1��mҹ<U5n�[�U	÷���Z�sV�M���i�&R0ȯ���T}{��l|1�GFjd%dbn���k��|y��m�VF�I10����N��L`;�lf3�4}i��yp���Qu<��d���:ݷ�g?����h�7���n[E𙲒��X������!wYT�2�d�]�8ɗ^�����X�-6>~�XU˄Οr47Q�|�b�������M�a|�}r�S��W�l�~H�*Y!�P㣏�q-y87�![���]@ȼ��k��c����ǛC>y�ɣZi���0�^z�$��t����\G�OR!�����lD[l�,@���]'o$?e������a�CI-���,_~5��c��k�ſ)�X����#Be�\½?7��Ed(J�\
Ւ��L���c�Ė{�U��"/�Cм�d��hn��ia�4E���
?�EH��k?'�O��L�g����S�/WNZˉ�����6-V	]v:�Gd�<-�j��D̯��R�|�4�g��/��C0�c=�	<1��"��~�˧���#�֦KȻ������0K�X�]���(]-tI0�{>Yh~8+�c���0�a�{.��{��t�v>��I�7�����u���Y��"�m������Q��42��9�V#cWz)���=͝�w�w��{������ Q=V,�D{��u"28����������G$2���ru$`�(P���]��������\Yk�ZWTR^�"[��E�n�.^f����s�G�0�nHy�%��߀�޼������V�Z��(��j�Bv�%���7a�`>n EZz�>`|o��3�{�m�Gي�IZ�� �ʀUk����IM��K���ݯڃgt?h`]MM���a��P^X��?�'����f�yxk���p�GoMl�We�'�������<���Kx���"A:��4�`��C����.�	]�������+��LCa��gZT��[�#�nB�?���u3K6�Y�{�&��!f�d[��O=f le���Ɋ��o�d��/	���2��k�-kq����bv֏�*K�B@�ZX}nw	:u�,��+��r��Iw�!�:5�B��T�H����w�k�
��'�!"ӴN3�-?3��M�A�cm��W�,���a�"j���{ vy���$lI��)G�۲7%��ߕ��<�e*����)4�r?�4ۼe�CH�|�6�?K�owvtg��A��X��_D�FD㿻�J��\�v��߅m$I�塐P��w�Q.�V�'��cD�74<ާ�2���Z���z����ET��| ��\(�E2/L9�@���W��
S��sLWK��M����M��:ޫ��Q�^]�6�5\����}#k:�9��oW�#����؋M0w�A��zSIЙ��D���V��st�M���6��8���\+h�l��/^�
C9k��]�u2`'�͸�?�r�O�%�jJ�����ph2@�/��^���u�y�NdY�|�L�BP�c��P��[`9ҭm���RT�<=Z��F�����+>��ce����iUT���鍌׵���E�<+�_9L%I�>�\�b�8
-����߮��/<���;+U �W[����@�q!aD�rCW��[֪z�����׫�Nv�k�Ga=��.��G��\��s�M�ݸ��.���9�V�$��p�,����K���1q
\������>�1vs�W�2T10�_����c�S�wR^F��i?��aQ|�v7���Ǘ8xZ� �����4��#S����S�4�,���Nr��Qa���{R�������#3��>�����hݐ�Vc_ �:	6��(#PJ yk�>aL��m��CE��Հ�T��|8"@��cK��	����i5@�%����1PZ&^�Aw��n��l最=���5���u�M�#��-�O�Y�S�	n�x�3;�� .��71�W9;A�?GA�l���$��m����9N'�8{K����AUx<�~���\dwg�,��qe6�sm��ucPJ��L��ރ�����s��ף��0B�q��d�(�{�M�( @Y�,������P��{��UoUDLBq��b���r=��۵��?2��&�%��Z��R�L"��?)�ǒ��PC���kg�$(&��^���!��:��\��@,�c¥e��*d�{�7@���t��0�E�!���)��k�iD���h�-<��$����_�2�rZCJ�����B��`,���{O��k�X (�����eWG���5�B�K���TC�