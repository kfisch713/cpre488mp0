XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����	� �d�%&#u�r� ���V #Sf��w����έ��4�"�t[v��"���ݍ��K����uǣ˒�n)�8΂W >�s�~T��M����1I@+g��>:4{<qҔ��c1���h_�Ac���ϧF������)/��v����i��7{��r�Q� ��������0&�x.�\� 񡊦A�D�,�i|�4|}!Ο$?N�}̙`ɩ��9�.�ZO���3��pTr�����}h�������D/�����
t��S��k;mw�(�>��eLCx>��6c<�@!CIKa��m�~鞽�E+):�ll�܅�UFr��4�ĠP��@u�ʞ
|1�d�ޓ��{���A�.�5�)�2�¹�[m�� C:aݕ�R��=y�K��"|{���н�����@,W�[sIm��vxY���ԗ^N��끑����q��j��,��_��%�[(��m�l�� &@�
s�H�F�J��Pݻ����=��>P�?B����D��U?��'-���m�����a,�ݴ�#�[��*A$f��a�oQy(�@H$�<E� �U�V��i~��/^�	1�a���:�7��%Q�(��p2�w����1v�q�v�4������%��'�I�P2UX"�ߏ���}F�*�����~N{��}qܹ�y�؞�_MW�ث6���I@�}�M!�n��n���޹�;^_����
��.H�l��Ʈ��czH-���a��%Kir�����XlxVHYEB    6346    1790S����C�>�bw�'t�����>��eX���8'�H�4�Gv�n����$���e���5�]k�u�c���${{@
����� �#�M���ΧɄ�f�dG��(|z�#b��Y�G	CY��qփ��� �
F�����H ��).��R�y��*����+�4^��F�?W�d��e�������2xCq��ǲ�`IF	V�}�i��Wsq%f�-�ք����O�	���q�%�����s(DD��J��#h�R�D��O�M�x5vL�=Kd�'�\Y�
�Ώ�:թ�u�Y%~A�q�\�D�YQ-�o���gU�����O܄�l�dژe�
jn��徜ɹj�u�����
®�.�]1N��,������b%�AUoufI�~>U��W)X��k7Z)Ȉ�#Fp�������xl^���+a�N�{º�`�'��+��м��$��2�z�m��U�vͧ�~�&��kuxP�F�IP!A�$�}�n+�Y��̝���I>��*"`�*��{��� y��s��W�o�,���(���uǐ��=�]�3��X��B�	�6ip<����LJ�ſ��($=<�r�}T�������b��lO�m�B�{V d�P�b����G���A��:��x���q`��j?�W\���؝��!�;�C����K�,�?w?Ȃ#����vcN��p�v�Wͮ�LԚl���������;��kp�1P��Ci�1��6�IM�,�o��m"f�-ϔ�2٣(i�/|��-�aDƫ�Z'^p�	�Fw��	8�mPS���O��&��r��8�S�̸�*+8��x�\�@j���Y(�>�M��E)K��M�{��$H�n�r�Kf���\o'�k)r��?��+�Xӻy��UC_���`���1;T�+ij�70���P2��6�9f��1�$:���dN����ы>�\Δ��a�b[�=�v� `��bһԾ5�"����.QN�cs-u{�ob��,���b����;���Ά����:r�X�	��>�:����VL�#`�
2r�^���͙)7�׳�	{�)�?Y5��q�0�G7�?���C>����XM�M��8?�����`�k��l�gz�K��=��!"N����?������Ӎ����b�t��Y��`�e񲻩L�9�ڰ3��rK�����B^a�;�5��'���z�lܤN�Y���sa��x=��J���h���@t$@6#���h<�v�{/��@RR�`��F`RH�(TZY�k]Q�>��1�+��Kk;M©���g����ߘ�ײ�ݩ�Rj�Ūg�O�+�V��'�	�F�s"�Tf2�0<�h�lH����
�g�'����r�~K_S��?l��x�ۡ5;��lu��,���.�T�t4�]� �kCgH��< �ry��/��`^��j�z�=d�Ɔ�[�����eQw�����#y���L����x�#���W���2~�`Q��ZW�h��n3�{�8��8P̠h��kIs"Nì�Ml<k�};���;Y���Ne������RC��^Xr����/�:kHޢ�4 ����B�m��uMELl�p��-)���k���LM2��C��=�ZP��"�W�#�������H7><ԥq�ū���}�Q�Q5׋�v�Q���[���6`�M$��Pd��� �#�!����4�����ʙ���ʱ	���~ߑ	�F�F2c�oՆ&g����9[�����ʍ{�d'���2�U�*>�̍	!��1��R�X�S�a�\���.�(P�~��ی4�&�v�l@NQ��J03$g��������K�6,��܃��]�z���+'4M]�|d��F]��߄��HV�?��P�Z~�C�h�Z� X�,y�ެ�%c�pV/?j�a�ٗjr��k��*a�����q������6V����75Ѳ�Au:u� E'��HZ�eu�w��8B�0ٰ^�'so��㤃�r��E6,`��G������gY+� ���%
j�U��}~�	����5X�X����+g-0�<�^m���o�u�gN��@4.��|�\^>�2�s�n���ng̷B���JIT��2Td����D�p?����9=����6aX��&�g=
B��q��x�����,'��v�Z֫���8|��3�d�d�M���S�ы[��eV�o$�,;Eq����#�ʬ����N�_�;&�4����O�4�����u�����;����*h2��uc�_��s}3� xDW�k��'�=�����!���#؍�K��ݥA��tf�(�ڴYde�-�@�K���Qœ�"='��X���N��I���MT����7< ���^���Q�ܸ������I��$�!F��5�}	F�Y}��Ur����Lr�-���t<��O��Q��|tX� M'"LY��[@/�-�:4Vk��;������=�H�x�4  y9d�����K����勱~�=x��S_ I[P0>���E�+�F�9I�i�F��8o��hb~�
+�Īڭ7������W��S���8mX�;~Hi�\R� ��������ԇm)ȰBi��.�&@��M���Nc��e���^�����@L��n�s�S�Z��7����1&D�)L�|��N"�0�>$��A�H9Ov��	~���)���YM7l��f�Eu����78��n�/̇�^*�ԟ6��8��2֟��x�k׎�?�%�N 3��?3[uS���-�P���h#��Vi#!i���e'�{��"b(U[U ��
�5�),y9x�p�r���V�)_:�4ىb*�1��_���oj
Ϝ�� I�������}��d����2v�����.X���Fgx�t��VX�	n�eW�-���8(2�%��P��.�'��p:p@n�p@��������$�/>���C��+�@h��a����ɏ@C)ˉ��q�����{��6Ě�8�;��21f���������]�Gچ.�.��<�n{[�.���ڋMр:(ܷY�4!k�`�oay+���2IE���2d�^VYl��M�|omfp��w����k# ������������e[M����ٗ��sy7/m�p!wg(1� �^>�#QLF����B���"v���izƒt,�	Q���V>��J
��lwأ�V-��{�B�n���"�_�F�#�ɮ��~y��p�|��Z���Z� _��
g��ưy~���/���o�[jT��m�}��Fr�8&�S��F��^���55�	���d�@�\�(�I)��i�dW��A�����hF�/vo"Kq�V��S"��;cv�b�K� !�c���"(�����<�Lهu�a^|�E�4���)�w��=ɴ�Ŝ�-j1�a� �V'pq�Q+�����_oh�S���-Hw�_�9_���PxuG?�.����@����o]����,o�J����3��8Zq��8�ݵ�V���[A�_q�/����'ԑڴ��������kaN��F�¦�j�0CZt�Pw�оfC�J��j �ky���i�+��ur�P=��O�oǩ��,qn1w�:|oC
5w��\�<G.�Dn���c��Ϭ`�*Aۅ�J� ��+�8�O�'dyw���%�*�~�]3�$|f�B�[��t��bM_<s��j�C�L� �4�������jU��i�6�g����*�3�@�hGv��+�\W�5e�a?)CT�)�V
Ο$�R�ʍM��8ɻO
VOW����V�	�n�x�E:�1����/����+`}����'X�-ڄ�#��L#l����ooLVYB�G�K�-l^*;V�̈́�Euzu܅)��qB|�k�{�Ǖ3,m���w�܋_�b��~r��(�ɯs�<E�t�/}V�[�n����bIp��%���|'�g�f���FsI����H�i���Y��J�p����[�.���8�������xiD�ܶB�s�{����P�X�.��C�׃�S����d�g�'���o+l�����v1�>4Ķ�wF5�O*�f�> 7�,F _ ��F$Z��6����<NL�a�m=h>�^�k�s��C>Uk6{������!�M+�I���b��+EG���-{?�h�MO1����I��!5,Nȳݹ&.yF;C�����/J�PY�>��Q-!c��6V���n�ڑmVL"�����(H���w M+�z%�69�~[E�TwB]³�}����^��7����Wv/VڑX�'�dE���D���D���D(�M����F��)r�nd��"B��v��c�	�ZٿoۊkE*g���*K�V��������F��E8CH��B�h�V��O<�mP�VDC��U7��\��,��#ȓ˭����m�D�M�#�(���]0��Ҥ�*����#���bM�t����e��a�u�,����&ƫs����z�[5*�V�p6`?Z��hcZ�N�����RnB�{~Tk|���x
&�w�m�C�U�g.�4L���fX��6E�+>������6hS� Gjb�z7���UAw/c�w��9�t|!ԡ�R���f�pPa�W��� �dSHw�&���V�N3��;�i�uma��z�CZ܇TPF%6w��%j���Fs.�jty	�JG!j�2H�_ w,0�6����
��6��۬Q�-#��=�m���lA����K'n���>��yj�Wl�-�i�E�_��jɐAX��0�ү�^7,G'�� �H�Jeq*_z
�%���m�l� v��f�Wa��~;nM�.���� ����u�;+�3�:����DGJ�>�*S����fv|��*Z|���^�ʨ�����a/�Ћ���q���a�O�r�A��h%Q�'�-����������p���PF��S�����0���AZp���{œ�MGb��?/�I��K���k&��'h
��~M17e6|Rf
Wft@*�@�[v3Q��
��*qEn7\�B��f�?�Y�Ne(�<a:��?&�mD��:i�IA�^��|�::���1�I��#��o���N��窧��^e@�">�>��@�SZݫ��G=E-��ʂ���υ�$R��R�2�0�	gދXM���"�<c�O�0���������?ih�nᡕd}b�1вQ~"�i���Vź��Q]�'�_�u��L|���[/:֕��yF	V�A�ȒʟV����1�jaHI�+Ć���EO(�5ã��d�NE�hm(��Ťt��\���y2>mz��,��>��q��Q�򙅋�,~��0
P3+5��e*՞S�`4��G��^<��@�쐥9kt���v��M��#~s��[��j��I���1!I��7C�n��O���/����0s�uhY���̝����"#w�%k�UR<p1j�&ͱL��:��E��fe�^L�|t]U�-�n�2;�4����z��c,|c<
����Q�g���ɛ4�ɠ/p>�EK$,����J�nǇq:����0���3�Q�@�|!L��vE-�g��rqTD`V��Q5�68�N̯.� *�.�&�\c�ku�'���m��|K��LC��� �D�U۴��41I2́��ͻ��0Yv�$�j��&d�e��.;p���9{�B��;&u��J$tfX��LxE��1��ʿ���3V���P>��Bi�ʖ-PǏ &�����G@J�~B��s��$X%?k	�� [��/[��?^�P�V(���%�842���t��2O3��rM>�������7g�lo��6ω�4e���6�1�6�l�A��ܿ.�,��}��c�E-�³j�s�0��r߾��;rL�U&�>m�`+���O�g�2V� ..k��ʣ)��l2��na㦱?P6pB�0�*g[:�ګO
��Q�6�� ��Ŋ�<#��1�zK����bb�͌�