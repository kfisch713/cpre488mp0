XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���0�jl�VXCJ��j���bڪ�[qL���d a�	�h4���#L��U�V���+� AO�r���:���p#�>���]���
I4}>�<���ό=90OfS&���Fr+�&q��M��h����{�j�5�0�tn%��M��=��5A�����71�n��J��`v'G/YdY��&V+ƽv�`�9�ޣ�9�a�>�.���*c7d5Re��c���5^0�{mI�b�.w���G��˚ƕqm]|��(Ƞ�
���|p�����j�ۆ��\8��]��l��wz�/�
���h<=�J�3)o�~n�bp0�ܵ)���B�G�Y�\�����8c�q��pA�ݛr���<�6��7S0{QZ�o��O��)�#[˭w��@n��1�X��7��p�z�X��eH� �a�-�{�8o�-n�I#dߺ��I+}���PB�C�x��q����ľ�?���(���6e�w�Fa���*��54�E�	^+�e�G\�}�H��d&�d�tD���Xa���>"��g.ha�������^Qp�m�.���&s���B�������1	�|m��F�!@*ڕ�{5�C�p'v�V�c7�Q���q��#�M�"Onm��(|�4�퉞�$_*�e��xV�����MPE�D�n���ĳh�ZU6ǖ֫���ZƂyg{�E���U�+�U�HF2�7��I�9."�O������DD�� ��h���;G��b���`ln�g4�q��e�	��K�*�K����2-XlxVHYEB    1853     810�*o�>��]�]L����d�L��{5J�e�0Dt�"����������Xl�m���9�|��qJ ��{.Ű�/�|Xv:U�M�Mp��u��������/�j%�$��r����N`Cb8���E( ��$b(�D$=��3e�wtY��*�Y
D�����P?�?J�Lѥk��C@>a�؁'v�q����6�Hu��j+x�<!ϰ�-�ZW�'{����C��G�����Ç�0(��5Μ�ZA���qMSd�U�
v���iS�ߪ�o��c��KX��uBM��W��/�ٽb�T�[�/��.�v��jcy҃�7�1ڼ02Й�@m���z=J����#`�=qy ��W�VHm>���������{-о*!W�)�KR�12هUr�n�K������!V���Jo�}����ef��+�D���\��R�����ё*��q����q�( pDB��R��˅z;Ma���]Q�tE9�dĳj.k�:^VW�'r�ª<r��ll��fESy�C��+N5�9f��ך�χ\���BjY5��׻R���������	x��M"ǐ��^����Ug�.�j�>yj�*�#5�B,M�D��ٸ�'��PkY��8��-��s�����P��-�6�^�(�a=t������
�n~�&��[��q�خ���s~S��v%p��d�� �Q���N
;O�,�/�u�r�'U�ȹZn��I�f�)u���@�`������)��a�&��"���"$u�LŪ��1��s��A��T���q���7�`�1.۽s�%���c�rQg�*L�g�.̃�J�p�G���n�P�eho�c�}���/��x����o	<��+�,+�W���xo.�6��������}c�Ԍ|]���P�'�#m�d�̗��T�d� �^�-WX:�\�!'���5۰���I�	&B�#6c�lM��9��Yv:��k֚�iAg[�l��Y=3*|$'�-ygC>�#uC�k��TT��6"������Լ��]�/�e���k��gS61uG��i���ЩJD�ui�j�_H��%3S�2+7^�6�F�)oG��+o!�s;����LjV�hV;�� l蚎�J��=�� oM�
�S�9���*�ޱ�s&��r�p�<�����벒� �}7a��F|8 %C����n��Vʐ27�;� <(���f]�ڄ+a�9ڭ[��N�G�n��늒�
�L�Y�L�V���%q~:;W$rN=�S�2ou�Ȫ9����dxp���5�ku����j[��#��uz0۽�n;�g�d�w��h��^Yr�x�}���{�6n<�-ք���؂�),��w�m����g�P�:��:v����spgK��i����L��]ƍJw�؝D4=c�GQ$�$�xT���9F�ty�C�'1��ٌl�?��Al�l��w�ii�Y�۩Υ58�?�G�.f6a���t{q���On��^��)�J;9�G�J�n�����	�����5�W���T����-�s�1��W�����Ϸ�m���m������BzI5"�y��C.�dp��~�ᇾ9FE%���
��-Y1��5I�	����C��ۥ���	�����)%�F,C0���&G�t�]���BM�%�(>S�;Q[m�����dd{��wa��Cs�E�mD�B�VBm���i�ׇ^� s�*uN=�G�9�F�R��Aӑ(��!r'�.M�w����Mp����ZB�}r���bg�ז�ɂL��gl��}H^��_n�_oTqk����r�s���y�E���9���P��R�sr	W�'~��`����1��ݨ��wԀ�S�܂
�f��ͥ�����鵽���$�G/V5IK4 ����l�6�w��H����9Ç�e闫5�Z�2q�|�&T'B�����������	{i�F�L�zWN����A� r��ǆ5cy�TR
m�5A>��ҒzUtG(��X�=y'�ШR�h�H��9xه,>�M)h��pܳ	=�m�e�� C�u�Ji�{����