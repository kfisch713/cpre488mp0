XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��fgi��E���\�Lz6�z!H�z �O�K�X�~`%��=&�����l��i0-	?��7�,%�n��r<�f�F\���j�^��O�p�cq � �� ��e;��4��+h-2�T�@���pVau|����r�� �3��~Ov��|�MɱH��-�����0e:�3*���C_2�R��]Z�1yѩY��ʀS��\&�.J��PD?B��#Z��J�It�*��TJ��$_����a�=�]S�+ �U�F�JZ�5YG���m@'xrm&�)�Bc�2�2'�����'�レy�B�gs!Js�}h�p�ZGFգg��̢E>��k?��E��!J����㝥��T�JR$s#]�g�,��I�D�1�4�o��!��b*�I��S-[_Dx�is[k��i�/P�܏]���K�&|��ڈ�(ToN���Ţ �M-�ï��R�_���ͳ��M��e�.��D8a]V��gO�)�#���� 9�������N�b�9tpS��_\���	c���~Cو	�9��ŏ���Jt�Hk��uQ��J8��#�Wz����ߌ���#a���7�}�*i7�%t�Ov% 议�-�s��T��?�g�h��{�'��S#lPQ(�%L��2���<��H���V[���pn<��
����i����A���b]��z�b?Z��iR�����A|ǷB�Q���Y}4��l�nb�2����?ʐ,vC�D(\�+�EKk�1��ᛨ`�s�7R����)b x���XlxVHYEB    3fdc    1160+E�!�|��Tɞ�D 6?�<����d�wi*��5j|�sK�o���r�Ѽ���mɘn�˺�����.�xm#n����5b��1_;J�*۬�ؤ��6X�����,�v�&&)xnԬ��ȶ&��v��ބ8�ߟ.����+{�"�>��9Qcy����f�o�%��p-�\4"�s��7���r����ֽ]{.��!i���\��gw{; �b�x��(�}�m�1�C�P��܌Ľ����&y���e��/L4��T4�����{.��h��O	P6Pۡ�tԦ!R�g�C�ϨHg��0*e+Q�訙���@� �r#`���/���=��H� �bc�#kă��C�����!�O�V���=g�1��th�@��a�>%�فC�l��E���t�8 %�;۲@x�:��C@W4����C� �O,�ą1Ď��Y�>G�@�;%`*+ӊ�þEE��c${4h�R��X{����~-��7]a5��t��D<�,5���Gf����e�D%�%������$����U��{���1G�$����W�Ǥ�O)�I(L������H/�jJ�6]E.�գ16e9S$��z�B���.��CJ�=�W=[�HLǟk7�+i�K���+z���ʱ\)_ɚ����?����5h��'`"o蛵t����\��p�_����w�y?�B*�]�x\�B�PH�p�ӭ<䟾,�m*Z�E@k=_co&[Z&�C�)��Ҙc#��Ұ�~%=+r�q�i,/�'ޘ��W�ߋ]���/�)tQ6������+ %��".0� C�i_M$T^k�9��G
6C�F��dl�h���I�����䶘���T���U&�m�
�O��5�|�1֒1y`��1��}��
ew�6�q �,!�Ƈ���-���b�d�њ�0�c;M��Ԃɾm��\��S<�l��Z�B��j���E����`����[U�Ɗ�ͬ�l�	!Q������Kc fm���A��<��ܚF�p��#��47eXM�Ղ�6��
��Y��c}�����۸�ÙrCr�l �v.h���K����~�$	id����Ύ9DMÍ��ۨe���]J�T�s	��F���D��u>�O������ҭ�LP�e�%���������]\(��)�k�����xX�ê��ܰ�;G�����"墻u�,�S9��x�L�MC{�m_IP+�;E�b�y���j�\Ľ�E�_� ���Y�B ��-�-���[����(;�!z��W��T�eI��d�J@m�:"$a��z���}���;�QI�^��)^�s���o'�y����8\RvS��|��d?g:%P�C��Yx^(���ǖeyL�j�^ZH���;ޓw|��VB��w8�eG����y�]�;�ҝV��D��a�[�31˵�-��q-|���W�_;-�ؐs��p���
5P��<�.L5w/\թj�5��t�\��
*W/���Νl7LF(?_�V�^6�k���t��/�3�u�M��s}k�B����R.�; �C򗾟�HKs�T�^wyZ	0e���Y��i\з�B!���¯�і�5ч�'x�a�<g	����6�}ƀ�Z��:�o���i[-G%b�tL7̴Uϔ���cKOয��5B��⍓��P;����Mi���	G���w�$��C���🷼&gY����� ����ݡ�a�R�`g6�+x�>z��;��|!�t��Y��b�}����j�u��Ԕ'.]�:Փ	)�Gg$QVH�t���GN�������6���첓M���}:�!֔n����+R�Np�q�xL�Xc�U�O��p!�d�q�
���%���W�{�CI�5�BM���	���@�����w�u;%�<a�|A]����鑽P����	�6Nd1s�Μbn9ede2������N��Mu��B�^֏S.LU�\c8Oc������DP�?���I�th��H�.�Qӓ�)iL%�1�Ihwp�PbIQk,�a�,���.��x[*���ڱ�z ��)L�����0q��o!i'��x�����8�`	F ?�_q���5iҊo:@5��Ţ�9
m[/��v��G��_Ie&0�H5p+��3zk@O��B���0���~�'~w;<H�p)w���Է=������6|Z�F��sKݡ/�5){�ވ�O��h*I	_�����n��d���F����) � E�m��f�%:�R@w\Ǳ�Ϟ0­�RŖt��\
a�G����(�R�{}2�mD��b9S�fX�N�u"RY�*����Bۺ،��F��b� Lw%����)+�r��h((��}��q�/Q� �������Q�<tJ4�ح�݌�i�U��]Rv'�b|ps+��C Q8�Qi�\�=Z��x�R?�"�x��l��7#�2(jy?��9������i��X�g��~b�:\~�6	F�k�^���z�Wyt�K�I�Yk�{���4�2U���~d �vn-��M۱�~�;GZ�3����K�\��i� �Ѳa�t�_���#'��dED�N�"z��|�4e3�Av�F����n}%�������(Z��]~	b�뮍�K7.�s�3�a<9�2�H�|3b��i|5�y]��-��Fj��j$ ��&��}����G"��g\��
㊫�&�����F �,��7��3o]����܇o����]N� l�H6	Z٢��A���6�ʔ���и�g�$�xa���wL�a8sp���^W,2[�r��vU�+Y��4�����+�P��Q���� ����ݳ.���~�o#��NM@������5�d*:o�5(���X�pApW�P|��B{e�W+�7y�!���� ��fm��,�eA1��?�[�8�؇ڣ^C��`))]~�@}��}����7]o�lw󴸮O�['�SK����=��'�=$ϐ��n��p0x�����IW�1�'�^=��FV�����Z/L���XҨb��*sdH&�k�J,g���%��6ub��RheF7��c���Hں�VYa��������ý���?�^vK��b�̏@�75/����Q��NFb*c��p�W鱲O�S�ϒ0���V�zeq2�9J���Iy�N�0��D��:�{s�v�l'V��Zj!�֜%]�^J�y6�˖u^�?$�d�5g�o��<��SC�:3�ȯ��4�dy.aO䐊�԰��aR͉Ĳ�g^�h�:�A?#��0E���W�	~�l�v��5h< ����iB'w�Z}��$���4�f�"5ϨD��W&�HN��p��9��e�:��yji�uz�"��m��"��?�0~�D���� ;� y���m~ё�@wI�73����$�3]Q��Hha�>⧺}{n��
��Xg1�r��~|��ڢ��Ư`����'r��VY&��Yv#8��a|}�4Rwo�c��5GV�����M4<_�:ى�$C7"�H��5�y6���A�ʚ=O���9��	�>�M�c�c�țd�C�&
�6�,���@gĤ`N��t��<E9�G��d�2�ZdPU���W(�W�
�p��<L�)Kď����@��!�x�笲r3�9�����Ⲟ����4��I�5�4*҅�K�Ǘ���C������&��fC5I�&���$h?�8A&�|���)�ȚG��[��o�,u�و��p%����!.O�p4zܨ�b�Wȳ/��E4�Ȁ`�����+r�rA���O0��sw�Y=������"B�T�Ep(���$��Q�w4rӵ���+�ҟ��13~PFZ�n8)��5��\I���#�#�����p)��j;>W�jx#]L/�3=r��b�m;k�Ӵ�$븖�86��)�m��'���;l�yOQ�F���Lȯ6͔�"/H,�����-����<%��w��0�Q8<)�(� j ��Ə�f�FE[	�u�0{�~ߜ���L���[�Ǐ��,k�+��-�!o�4q�ݼlJvs���� ��g]�Q�[�Y��O�)HV�e��u|]��6��3��	�3��{Z���	0�*�E�?�$�s~7�����lw���1��A�����ŕ.�����g��+Mb��{��<�N�X9&������U�<����؉��<(�߿u�Ԭ�]�����,$ [�p,����e�CmDmz���$���CO���N:�nN8�z�����=��MO��|��?���<�'�2�� �}��m��IkL{��5�T
����*��~O+f�������p4����$�8F0�vxu�v�h�vߔt�È@�U��X3Ƽ�u	{'j��3J�}�əH��� ���/�1"擵�n�n�������h�$�UQK������E�C#�V