XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����'�O�m$�_{D4�!�"p/b�y���J�|��*��$i��<����ڹ���I�x��iA�e4���ÅG*����}eۼH\� ��I�m2�_-��](yS��Au�0��#��>Ԉa(
�>}xĬB�w�~@����gCm��:g��|�r�����.\��#{�}<�O#�n��H@8</��&kQ@�+��E^X�V��59e������C��@<�;#�������:���Z�bu��bD�β��i}P��C�x��ȩ�<ݚ�]	bԵ��靕S�c���̿�H��D����37���1d�iHa��RE�sp)7 S�E�����ر+R�SI�6�=E4I�w���^�>H{_�iܡ׮p��픎�����5es�h�1@Ӹ���i���(��/�p̝�#[����nB�%�;�2��6 	��5�N����0Z���������G4��;c/����pӄn(�C��E+�,V9}� -4�:��#��FH�.q=*����2ӧ.��@���E�dӓ������S�*)�A CJ�?���}K���(1�~�Vx���V�q{c�Ui��(	�o�!88S���t?Ör@���L�tN�K �~�Y�2���D�/���9����]�̆�%-�eڮ�9xC�n��*���/�\�쳫{��2��6%��z���1n�a��I^���2ǌ����uv�C^��5��lB���b�6�Ɍg�� �&}��1&�vL�)��p����jp+U��X��l9�d����=v#"XlxVHYEB    3fdc    1160',3��Ǒ�x�����]_�����9�a3�k�+٣�^���;"`�e����0?S?�:��ܞK5����p-7�����eR�����?���82=X ��k G��5б~)��cxU)l`;1^��m��4'��V:Qт'��§j�N躊��W��i��n�YS��h�	�
�?���=�н'
<��]R�a�����k������O2R�)�hҸ2)�޹M�B\=͞��o���U��o��e��Q>M$���!���O�~�8�j
��������{�	�ex!��BY��e莾�>���0�h3PI�V��s����{�R��ɀ'�F���d��+`e.��D#������Z�n��Л=��a&lw�M<N�H��5��!�ٓ6]֍m3���2��=GI!�<�p�#�k4=I�H��F3�r�o�@��	ƅ��^7<��ag��L���^�=�I<!�P��p{a��U���P�����Wa��؈��m�Rѳ{#�^O��ZX�7��Fr5>��?��q�-�ڑ��8O�����!L��[}�Y�+�~�d�F��l�n�Eda�+�+��z�rޘ��Oi[Y���^�S|�,�ݼ�vr�X�
��� \Z�>��	�#�+i�/\��U0���i|z�y������pjf���M��ǃn<�;E; W<���Ҭ���Ʊ�-���/2�sF����V'�>o�u�lcSA�Ac�=l`FD��ƥ��+]���u�Ls6������u(n���"���8󾰓��Jp�yD�X)�N�NO�멻�	{B�hz3I}�?D�E8 �?�" �`k{߱@��GA��r�p �^*ظ�4hp�����A{���hV���V|M"�t�y��}F�z�`��M��0��)P���l�>o�'�D@�߹�1{
(:���M1�0�����?�tE��Z������m4r�����s�w�con�B���ď*��<��
�-t�f�hcO=�cGM�4����0��ȵ�5� x��lj�o�sX���(޵��Ś�-0R�=W�J��k�PPU��+�5��~W[��P��+#h��YY��Fqa����Ø���fR���Ź�5��2�"��ͧ����f-($�(_�HN�l82���c�:m�+�;��S]¿vG�bhǚ�S�r�&>�w����Եa��Y m�Ld��@���%�$������Zn�-@ ȍ�<A5�������`yܲ$Ѕ���2�+[�.Ab�5�p�[�`l!7��5�w� D50f�یsޅ�P���ly�~�c2��1���ڢ~?��B�H��� ��?p+���j��f��P[:�^֝�CЇ�1����8��@�rt��bU��n���p{ޖ\z��ֵ��U'e����/``��-9U�� VŔUk�ah3�:��V��`��e�Z1�e�O�b��K��r0���aj}�rH��i��ʳ/~��5��*�|����k� Y�-Nc��!�����]|NŻ�{ɖ�@��+��_@�!�S$�hH^��(z~��X�cеh�����ڿ0�4e�����*�c���B��'�.4|�|��ws��(J�
M��i���3���!{M�KYĐke��7[��;J��o�j�~�\=؏�j�ǧ�iT����i)�"u�w`g-�p��7�'��+Ŕ����o�i�p�R�H&�8M�W>�>A�un;�S��y�����`c�H��a�r�.�9��LH2�2�J	��<�}�dH���,����[�_A	2������F��h�X������ߡ27�˝��)A���O��޾#�,+LȊ��R��ғ�����7e�1���b@�	GY7��H�ᑶ�W�	dz�wA=��v�}������S-�]��=%�1JP߀x���j[r|߲�&�!றoG���`����`��L���0 ��(	���=�ۊ��w���t�2��+/n�����*��Tz�dS����֖3ص��xS:s�;�L���ypHIÀ(+��^�FFG�+�3��E ��[��j��.�[�"�)p��o揂dR��W]��-v4W���
o�#7�_���.����*�	����A��\^���#;��[f�����q\�r{�5�r^�i��"��|+w���V�dGdUp��B2e�8�}{6��T+v> �� �E%�#d�sjWq��	9�d�G���ZU=���PUQ����������%�2�lܪ�����qb�3_8K�6B����.akI�4X@�k�{_'�S���Oq8F�Ҿn4�e�8�B��xXS�N8!��2$� �J�u�N�d�ݔ���N�����4������vT����]���(1��HF;T�,���K�XL�Օq8Vo)ߟ�Hk���cxI��G8�NT�%߈���?ߠ�AyhA�z�X�d՛@~/��|u���:?��b���B�{������0�&):C�v��4U����O��J�җi��Ù��7�}5����ܷ����^G]�4]��0"l���%EBa���ܶ3��Z5�ܛ��K)����R�&K�Kr+��,����bt��:�&{���H�@~X혡����O"��q�J�s������J:J��.��P��|���{2��f�n�'�@8FdAz��se�
�5�f�a��"���wc�w
��,��Rt�I�v9Z���e��J�)$����{v�I�fM}`���|4��������y<�'����������s�tt�'{��$H�V���?�B11f�]�eZ�x��s�9Б���,��)'���8�}^/�!G
r�F�J�,s|
�)��9��t+�#(h1��M%�c=���U��\0x����l�:|��¾��*��`��������.�����!= '��=�2�r1ꓫ��A�4��e�K�yݼ�Eyv؞x�+q��z7��������(��u�o���P��+)�ٚ<>`m-%�ܔz������ LN�A
 0'qUL�����v�Jk�^�^�Ā�����]�o����j���A4V���e�_&#��}�"��c���'	kB�A�{S�k5�bb�S��n$Nv#�̍!U���s�U,r[=�Ҳa�a:��d�T^����}Y]��nF�."T�O��cWU@}�	*n��\�Ҭ0�L|��	a\'S�J{j�� �^��2�Ø�Z�f"3����c�R<�[ �S{���qR����Z�a�0.p�o��- i����22��n��8���!���f�^+�.��cJ9����W�d[��ݮ�dƤ��9����=g�!��Gs~W��a]*$ �4l�rqݪ�G9�	��)��n�E|.�j	i�&'ū���a�ʻ[mۻU���#��.B\��ޠҕ|��Mŕ����+����{�Ma��3֨s�f�=���0�/Ǵ�p4 M��p)��w�٘�v�%����0l��D��뭁���W4�z���Z�Q&�?�Lԟ�֚p��i�)J��D�o>����_-�����{_�\G�_�sѢ��[J`71���m��d\�������|�V�Nc�窐 �[yz�m�Ie��}�.�u�mgV`��	�u�s����t7�$i��OD%V���g��sY��nm��X4��q\!Qo��c*i�o�����,���!y�n%��֦�����W-���o½/��qVQt\冭U=����Oz@�Qj�g�P#����RR�):�&�Yͤ�d�+L�h,��AT��RH�?c��CC����=䳾�1�-.j����f�ǱI/�\�p>�����ÎZ�=� I�~���#Nd|崱��<�l4���&�������-��m(W���.d��j��;�?%�]�&�Q�l�g?�-`���Es<ob�G�>6��},��Slg~�	�E>n�Gf�M0u�3�ǿ���Q�
!�p��-ۺ�q�K\�lOl��8�:`y7��m �y��\��2Ew��Q�2���_	R|j�5G̨ī�/j��M�|�DOfܐ��  ��8�����r�Bm�m� �'*zf4��I���+� �G�t��7_BM���NnwM�8đ�ѣ��.��\)�&�t���USB���Cf�������V�DXb	���;��0����m�	�O[ONG�c#HT-JFAf���1�!z#I�"��2�a�������l�}����Yz
7j�&�?�w�`��a��^R<�����4�䚲Fc	���QXׅ�87�45�ޝ�3S.��l�*7����v:ВQH醄�b�S5����K�2�XyU����/���xJp�¹/�"i��! ��<��i�ğ�m��'c�K��^c�xn��s����m�J!���,��