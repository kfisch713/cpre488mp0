XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���+�����:+A²}r��Ľ�2�vQ���iz[����IC�ǚ�I�5T 2%�>+�t�`���a��+1�������٩��8f�.��\h�1;Y�F�,���y߷�/8���+V�m����[�DU��c7�q�!�.P$�Q���!mK�j�b���i�+�ܠ yIE3w�4ð��%M����K��@�Y��h	<�q6r�F�}8O,N~�`�셜��[�Q C }�����Ý�4�u��S�(1��B,F e��0��ō��*�?Q��>����B�r��N6Z�92�����J:�0�!�2�̭�<x��} �3�ф��d�8�b�@�S�u�~%��.����W+i�,<ؗ��Fc�1⌡а�ـZo��zRW�g�`z�"H �����}@uqx�+�}���1A#��!S8$��N�N��ۚ4S���O˓c��w���6!���o�I�X�qb�*lI�(e���+,}K��h��M���Ux�h�����������]� ���"�,Kdmߝn�r��`nQ�ц�B�_X�Y30�mJ���)ܜ���(c��zZj�!j�0|s�fp9�>#����	��?��CX�>r�u��ĕ����u]So���2ʿ���{#�������?�iF/�e��m"����;_^6�G��Z5��H�����g�~���޼��^:7B�.���IU柉.;��C���~0Tx�^t�uC�|��L���� t�p�<�XlxVHYEB    42ae    1110��+G�3�j��᭭T5��lD3�zS
<����j�չ�~����=%�V\�)����a!\0"jۢe�{��[,X+
�t�z�	��}���o��u�B�W�>"�n~��F���B`�H>���s_����$�F����ُ5����aG\s����h�ju$�8�鱻���ނT�(N��K��U�h�Ϙ�(��S���&b0��@_�(A��?@v5 H�*_��̺�@�5�0[[��}�8���FcC�Z�+$$���us3α�����։B��@ �C��k��g6&]TV����1T�׫p y���F�6�����l^h��b�9cs̾QlX�z亳�{Օ���~��i�:�{3��l�$����&�U�"!z�\�Ǽ�S�����"����b��N;9���$�� �A}9�G���|�p�?�2 �^��0%f�K<ZW�DM	T�"X�ݲ���dI���	����6�iA}b�T$x���X�5mP�_�BT69��j�2���m�1� �՚�'o#@GK?η����&fĽ�$���p�<�NC��$<��	�~� �BϚ��V�_CR�4��4�Ƒ�wu���&�����+XO\?���}����4ͬ�|z�E�߰�OF�@E���9���c��m-����hFxk�ŎZ�e���W�o0�3��۪]���Hþq��)N��;�d�?�������_�J5�-ǋ��bN@Ml@����<k��o���4Z_�y��;�پ��K��<�0`��A�d�Lɐȗ��`y{�%�|�`�n4e5e��r��7uf��c"�M��C夘p��3x[��1�����^���,cuk���3�z��&'i{^!��E
�4w�n���5�aHI쟛�D�������/-;�@C�hR� R��S�{P�'�`�4�x���Ag�ޡ=��?��Kb(<��R0<'�7I�C�d��ֽ���I���sY��2r�0�P��c�2ʹ6�FI�Q���
�����UuJ����%k�}7�7��O�덦�U>�9���[��$�s
q4uq��B�{���N�S��)Cg��A��;�?�n��M����2�������̱QΩ1�9|�a4V�$���6���@��V�( �I��?[	�WJ�
�y����a���\���>�|�]�� ���R}&�|�����z._vx�4i<r�f)|�L!�
1^�'�<m���_vX����:Z�T��mI���`��QA� �e1m癰��tH�󢤹�!����	f����ľ-�TC�x�{�%P�6=e~%�R_����a�����z�8ߦ�lơO�}Q���Ԩ��O��-!.�:���D����җ|�]�
C���̘8�XA����!���ݭ�?�����B�� u��>o�����1>֑
�0���K#�T6�K��/ES@K����Y�.P-�X��%�&<�`DR_A�����.��[E9��b��I��w~�X͏�a ��F�Y��G����r�f�k`��KUt��f�>��P�P��u�q�҆P��g�B8M�E�3,��_��E�yoX��B�k8�:O�צni�'q�cU޶f+��p.[4dԄ,r�2H����{�:"��T�R��B�ma�=ha98����L�[�B7�)�r�Ή�ʗ�܈�rn�
���յ�v�I9++W�/�^mD}�hl}팻�L_z2C��R��]�|��ũu马c���<7Zi�_(�f��[�?�a����bue�&Jj�ˢ�����z���Ｃɔ �'G�ш��/W;��@�wO��(bb��s������>�c�x$b�[ϙ*�m.S���^qR�C�lzL��B9	����gɼSͿL�����-�@�/�����Aą��R|�A+�T�L}E	=�D	���9���I+g�;H'�x=�.��X�7>���!�X��	R�}�T��}e.\����Ћ��\C�S�Ld��@�t�_��s���mQG,�)��!�MIX���I�$���4�}��)�e�R�D�[vx���[*����=�k�r�kMgQ~�	�n`�U�"
�J�.���&��kJ�:k�{r�X������B����(v�$qw��L�E]��d+^��9���n*E�ag-Yaw��?@�
Y)�#z֘�CM7��Ɇ#M!���V�j�\�DP�� <�>�t�H.G�J���FiPk'^����Z���V�����V?�[PV!��ς���s�a�d���k��[�&�F����j�� Y�D�9y��ml��LY���/Չ��È�������loY�pY��r����:	���=w6�uڄ�n��TX�_B��k�$)Dz5���o1h�K�ɲ�a�)_?���%E=l��64״�5�0�b4F��ĻhJW�YЕ��~��t���#Q���
�׉�n(�\�.�~A:lOj���r��;w�%�1�ܤ{e6�F��b�C\3]��,Feo9R�w���(՝�����@/�F�� Aa�_}5]��k��8��qʐ[*)���f5�L3���M�9ҝ�-��������GM�J%�'d)7�	�R�n��j�6�\g�oQjc=~_P)M�R@�h8��ո�Oa��k���W;�� ��ob�\�����.�/���z�[ckR"��s�׽����t1��Q���aj��p�+�����0�]c�2Z��.�r�z^E��˞FB��_e����j \�(x���;-l��� Bs�L|v�ˁ$6Ǜ���P�Vpl�Y+�Μq��4FUt�(��J���'�xU�
>w��	f �)t�tׄ˦d�l�Q@���t���vC"7#���*�ƷGx�!z6�Ψ:���n:jw��Yy|�D���]�xd�� S	U"?�ѝ�󃾯ڍNXG8MK��t$�gV�W���&�<�D�+ľ �_ϒ��AG9�N}�AE��c���n�+s4�8���qգ��)���qPƮv���XB�Y,'����ʹ����h�2�]X���z��_v�et�	��K�He����y&F�E��E�K���^����SN�������G�Ry��	:Ty�TK#`a/{��-�)��**�*�lO�{rkC ��M�S�31�B�BYfn0�2f��}�dL����0�\�S��9V�UFY�K̊�켷
�@��ùK��������D��N��;����Bp�EL��(�a����b]d��5�g�^ð��ݫX�+�D�Q�HTLaU΁EĠ��Q�mK�o�/a�����i) �Vs���gd�,�GږN�Ne𓞕�8�
��(��D`&�P�)mS.�n�0��$�H��Ә�*�% z,���)�z�g�)v&�S�'>�
�B�ھ�H)���R=�F��>�9�E5�ڇ��xP�R��C��B?�K���[�9��#�34�n1@�?����-�,
ֵY�\��I2��:��߁�Jsاf��/0��U)���E���]A7������m_��~�G	�ؚum�O�Nn6R}˩��?��iݴx��Ѝ�8	�f3�H����j��mP���~]h;���!�ֿx�K�>"����y�H>���D�	+�(|i��s����ʖө��Iu�0��iף�F�?)���☂	qn;��c|�,� j�i���J���V�s�������Q�'>a鸬��X)Tj�'�x2�p�qGqa���C���q1f`�<m���i�aS�hi�55@�˳m_\os���֡v�!����H�0*r����{�`�_�e�G&�V,�/�!�8&�4t�jp��˝ �=�P�ʸ��jl��oP��.hy�3~u�\p����pͷ���h�7�-�_�%֘�)�����Ĉ�ȕ�QJ�i*���R�
�#*���ּ؋��ք�D}��6�Qr���oX�k�J���W��8���a3D�cgl�G���S�IT�|��޸
V0���_Fs�N58מ�i<N�eо^�8�s��z�b$�l�hh���"4�zl�C��
�0�[9�_y3υ})�SH�2��1!Ew���Z��fK{�9���<L���g��ۨ2��ڏ��~�����I<���	28�|{��O�j�/H�Z�]�NxC���eO�vm���t����If�T��U�`Q��2Z�Z�M��!M����٫WG�'Nnse|�K��z�pҢ���_�I�=�c��՜�����<�P\fɬ����7����+���Df��r��0�ȿ6����q��Ȟ5�1�M��ARىq5����k�:5���ag�Pv��՘