XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Bx��i��**�{��� xt���U[4��SQ.�~V�mp#ͤY��j@� 
s6Z�jW�Ro>�o�ȱ��K���.�����)䜈�o�$L�� A�����t���C+f��)W'�Vr���h���,��3��<��~OC�m�p��27�2��od��`�Z��@`#��fb~*z��7�u�[�Ǽ�j�5�θyTY���%�j80I�x0L�η�UI��k���1�",�l��M}��~����n��G��Z]Q;����s #Km�H��
`K2��+3��E�i��p\+�Ї�:v��TL����*��01ΩuWS��O2������0$6v�o����ށ`E'L��We��6[����8���;�q;p5zg/����OM�G���1��a}P�=-�0d��{��㈭�%M�bg|U�:�2���&�����K��S����/89�f�T������<����*Z��#�n��k��5j'�$q�0�$Tz�����-*)�:�۵I�I�S%�������cH�1訽��ܦ����������?�$F	�=��˒[�<[��iX�BN]6�²'��K�B;�����e���=J��
{]�	���O�.<��3�-=m��.L�Xb�x|��ᩰ�
�Z�-�PS�H[pV��@� m1��������׫8C��	�mfhJ�$(�W�n*P�8Z�UCf�\��k�>V������_�T��l�(���6?���	h�� �mAcXlxVHYEB    3b09     f80�`��D�&K���灚��ʉTMk|�h&��E�7%:�C�eːը��p�}�a�?CU�ږ� ۸�-��CX�Od����RMg���*�a�`��>�[��y����:�rUӺk��k�j��/��3�v»�"C� I-�`�8A{��w��r�Ċ(��rͬX���4�Ɲ�p����D4��޶�����f�?4��������:�%�3�:R�*=a-1Y`,6S�'c: �i���� 2^�en�v�H�Nb@��CWk��c*{:��vo�	=���-�3��M�g:Fb\_���s$��9�=po����E2%�E^(Z��(�0�5��m�ǌ���|妛��X�q������Z]�/�5B�mv;���)
o�v���e���3;��])��0H~�n52� �Wݒ�o�^R
o[��d��.�3�i���l�g� �I�:�C��ԯb��@ f����:�*�؞,+lv(0�T4�N?'��p����_���j4��q�s��ӷ�Ҭy�i���
�9J5{A@�f�L˴�( �1B�f��"J��m0_��Kl7�P�N8��"�}�,� -5��/.�Jɏn�H��h�&�c0h7n{M@~uv���SC2`��&��,�R�w+�#i{�j���;ƪ�0�A��)a��4	ui�*�[���ݵ�Ʊa� �6�̲���/�+�b[`�z_}+#m��s�>��i{TO��v�3*E�wX��+���n�p���3/E:!K���v��@��"��O�Tw,h�J���G�{m��S���=��5x^�p�<�p��eY�Sm�5�f
;1݋�5�1އ����?L�,E��]J�B{��/�l�a���%>?�)����Q��KO��<�ܞy#/���;�^zx�br�@�xv�?V�d�����}���l��G�p�.pL�U��&+Q��W�-���%��F(���V�?��Y$�+Wzj�DQ���'���X���F�n��<h�q)��s�?�D��Œ-�U�E�7ب}wa&R�:ȓw瑨M3�߿�&�m=!� �L�l[�T��c�۾aR�:����Bzi����D*q�c���?M�D!X7���2RbI�Z��%��3=�h���[����s�$�� iaZj ���ыwc�� �.��da�+��A��/���(*���Q�~��K�hY�>�^<Z�U�gd������a�$�91Y���ta����Y�nHs	`(�/U�%�
��	�g����,K3����G<MQ�+g�5,SEٵ� ��r�3)E�62��1U�e��	�	���@4�\����ȳ�h��e�W*N���EDp]v �_j�n��Y�En�a�����gM�QB�j�N{��)����$�C�[�A.���Y���g6��Lj����B@#��p�C���{B�:,/�1���hC��9w']d��D��U�!ԍSf�*�"��Z�
���v��Z��pOoO��{���P�}��-�@����^�e�����x�&ؿ�8�D���{�XrR/�O���!�N@��0"�#>���5`�ڀK��a�$�)	��nZ}�i�Z��v$K�}ý��
�=*�+;���3h�k�V[�UJ��"E.�Ȁ�)�^�{�N��&�Ig��50�$�TX�2۵?�����;9�/O
?y ē
���a�n�l���N�I���"�E���g-�x��$�������!T��в&�~<�,�'�dtv؛�.�Y��RQ_Dy/9��.��d�6@^�?��Ż�l���`��}.�L7˪�pY=�M^�����2��앳հv��d���~��F*�ָ��D��B�
$g�����n�����T�L�2����Ҡ�^��E�7��=Fۄ�6�>�X;+Y���D]G��(b�m$��۳��%cG=��b��.�X�M�� �)&�ރ��*�9)8u�YE�v*��˰�<گ�z�8't\oU��=L����&���W���f�( �C�A��7#�6��H�42S'���e	��<�.��o���*����S��`��ႎS�
�&��U4[Q������/
]���	2K�j�-��}��V@T�dǽi��v��7oX@�ֵ��`���x`�.����K2e/&���@T�7�-J�#�`��5o�� P���W>_
]�ē�����]����;v��>�s��i�ы;��"��/��֖��� �����S�l�·���2@��ے�(��
R���j�!��ѕi��F��{SH��M�}�-anE!���˩���<�w��Xe�Q�y�T2�5�{��~��H�����dՔ�k���/�f�?�I&+��S��v�{Y7�ِE�j!O�@HA�nt�vm��XV�GGN<F�U�ӠNƍѶ�bN݅#4���E�Rl8�z��ݹ�{q�,��/�CU?��V������/��@�:F�ץr}�L1@%��q�� %]Pb V��W�hC����)�j?�u_���1�C�D��K�݈JMsB�J\id�&/��,V��~�%��H�i?a2��x7W)e�� �v�9��413Q��1�y��U��-
;	��vJ�;���[:]嚀�XE��9�B�B��`�����2FZ�ׄ�h���#.�4d��x�`��h-�Os�[u�'#��UCv7����\I�v����>c�gW�l�;s඄P T�$�|pj��҂�꺾"���!���m� ��R1[V7z#~���� mr�H����{��bh�B���F59H�q��HT�2C9�d"'�0n�����b��u�gH�A��:��0��g>�g�������ӇA��A�Gs��TF��j�~N��$�؉��$��=<Wd��8���۽��|� �\e�Y��==�=PP�?x֧�B���.F�K�i�,�3^�����ٙs���e]�����s�DY*����Z����ꋝ��M�;�yx4�~��/\,[t����ϼ4?�K�.�b�9�m�	
���`{�ZVm;"�u�*"�=mBX��Y�����J�J��#�_��:��E�����"Y���[!#�$�@_�3�-氄O�>L&�:��%�h�T�OU�q� ���b8Y�H#�6��;O7��H���8V;�b�N������ຩo�˹.�F d�Gav�� q�'�u��;��+�?��>n�����)��aJ�O�sR��66��D�>st��7�bT��� 3Ut8���%7�5��Bu,��2{���0�>'��z^�پ�*� ��Yӓ�Mj�TH��>�:�&gE8?�����KG���Y�� ��B�r�7��pw����<'��m��(�D�Q���XdB C2��C|�]%�D�D�%-�Ҋ�i(�>�2������cx4�*�p�1=(D��v��ٞ�Q�~�]�9+x�l�a>,�����QV 'v�-�,`��B�D�jLh�Ͱ��q�PV�mTvI����P��h�b[1y�/��fcFB��Ÿ��^��ђ��_���:�&Vk����h�e��|H������g{�[t������j�Q�X}�sT#��d��N ��n"{�����GvޅW�E֞d^R��s.|≴�n�MR�v9��b`��
����`�ʋ�w�����Ӱ��6䉋D
�|"�cԛ���x����_\~�@�<�*Q��y)�4n,mD�O�Qj��4������0�d���8Po�8�1�c�2��!���y�m+�A`�`��s������Id��_,�J�h�y��y>�bO'��T�^;��d&�F��M�i3k稽����;H�� ��S;�w��q}�"Ty����]J�5�MN`��ˑ�I)E2)��2v� ���L�!�M?m�KH5�M2�uW �z��$�RϬ�%=3�}RB�u��E]ϩA\�ߖPT��g����qA�V&�Pp�l