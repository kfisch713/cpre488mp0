XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Kx�����L��%^_5�3Y��m,��K\<��4E���� 1Wׁ����/'Q����`������TU��=��7\���,?�7�^h���_X��/F�;�gV�U]���yÉ^�MJ�q�-p��)�S��W�P;u�������3�"c7��u�X_��.�GE���»�{F��"���X�}E��%6{!���BQ\��/@��
I5<�k�[�'��'����PzB�
B76��~���3��t�	��4<�>���圫U���И�O{��%a�����Z��,'���̸"�9���D��Z��?��W����799�zk`J��ֿ+@��wH��C���XN�y4*���%I��}�O�-"���Aދ��4�h&o�}(�&\� �(g3�����\�h���EǙ�.��b�g���i?�����T^��$	7}SmL����J\Xh���-v:;)�P�O��Z21ѐ�,9�,����7�:�l�����o����{.�K�]�R�q��_Dۗ�I�x���NL ����Y"������Ⱦ���s���-����j��(�$�����#oo6�>�YaQ����o��f1	���D�l������~�i�ү�Q��ǋm��y��[2Y�o޻H���bf["tL[~�a?D�ʗ���G��A��� Bi(HƠs�ؘ㟵9�ʽ��^ND� �F0[+<��BDԟ&��pS�w^����(/2�ݓ�>�}�������(�`���^1��>�����_XlxVHYEB    42ae    1110�����ҊI���ÊP:�5'0&�� ��yTP�i�+�
�j��
 "����(�ǶřX�\���G���eC�4O^k~�c$Z�z��h��y�+Jt
��-��$�l��C<�U_�`[i�h�h�?/�;N?�3�Ydi�b��\K�@�~��?��}�TW����A�Fx&p��
�H5Z:����9^{��-��(Izk�VX�9�?�¥܄��GX�$Q����1���%dz�OX(i>�F��jLAn��5�F=����OYm}��^�����J�����J@��U��������,��Q��j2��	�
Ko��0��,G����'|rm���V��.	��I[�&���	 �K�.��E�w?�߉�����"�N�L���Q*n5��X�(�xLS[�e�[TڋD0�ީ�״��Qm��c���d��r���i�x�������c[�Y����#P���N��E��=x�f楡{q�����<�G	X�V�M���3�T�Қ�(ߐ];�sm�"lfH�Az�De���Z���H�g�<P�SZv �r��2tq{龧4�I�j�WQ�%�O���iYg;j���H��ޞ_u��Q���� C��v���X*E�Uu�� �W&7K� ����Ǧ�f��~�D�O�qb�'_�FkV���<љ�(ZxS��YL��~JY����W/��g[X�/Cv`�,	���ŮK�F��@T��gە�ܢK�)���n�~�O$�q�i���@f��?�#��e�W���F}�@8����ߒV�߷�Q�J1��c��g�]} fg�3)�@&������(�rޠ��F�]@���ݑ��$P)���Q\���E�2�
�(��H}�z�\�U��p�2�*#?Tz����i@|J&�[G�/Ǒ��r)N�R��s�$���i�/q��=_L��,����ZU?iD�P��q
�|�_�=�sWڡ$�s�p����cƬ.~rǡ��ـ�,�è�>p�K���h����0�C���Ua�����vS-̧�y&����}j��$���: �:�\z��05�ingEr����s;���$n�ք���Z-G�cnf?ը0�Ag�C5���S��¼I�����Yk�|��@�6���0�z��gL�J�"x7�YX($�!	��ɉ����({�X( ��E)��vE�e�rE�$>���?똮�'����ju-����N9!���{����]}ʕ�/��Ϩ��ףZ�?�.�/T}Ζ$�vi�wC�t	NU20�W2��w�[�Z����;wsnW9��+���$'�n�ة�Ώ��X8b����f�Ī��!5qj�`�W��)��~��v��M�L�C  ��e<�Z���U;*3���T]-C���������k�CD��oN�ʬ җ����|�=_�asNm�d�i
�+2!2E��@��s�Z�N|�{)�"Ul�W��ę�f���6��`I@z\��vk�FYǦ����<��,�ZH�{6�KTX�FT�E��D�x�Bp����ty�%���MN�����ܔ?%�ǲ���Ad�OE9��w���l� ��6�,�n�����qi�+�L��݅�Ѯr�Gg�J�4BP��=6��ba��"�6}@B)��c�((�a&�g�H'L.C�sM����?c��EJ��P��i���j���?�pK+�Ǿb��Y���m����x�L����JXr��,�ɩ¡xn�)w6����b=�؆5/�~o�h�[��B�9�ziG�G�9]ؙ5ޕ��`�؞yE�����z$0���;|��;K^.2�,�	��vG�cѝ�D�=⤐s`��bߌ������o��AwB���ח�G˩(��j�۴��lX�z>�ೄG��"����� P�b_E�e�-p��]B����F)�̤���P�̃��Z湇T�!�(�
H��&T�����W'e�g� �n�"�����b�|��@�Q��Wp�l@�������a��U���CB�G���Q��ˈk� 2P����D�uX��Ly������\�K7.�30�+�[�4�����������%6����2��F����=~1H���I>%�cX�x`��z�_��?27E�Y�ݢ��j�,6G"�_����&-s�˜r-�*��7�����g�z�<�x�'��5�.C�P�SA�pP-"�:�t9T��Fr�����]�Ç�#X�Gb�{�L�0��-��zqbD��,&Q��'���=P\�
����j�*?&<]*����PnDkU����m�Yy���lЂ��w�aFާ�!�}z�*3�F
+��9��u�K��.�1��m�o�����G�n"�������$͎~�,2b5�?R���f�0-��e]��?tr+jY����a�O,Zh��o�F�ܵ��~�OY�%�\~/~&&Y,�K�ݳw	�+��h�kZ�dtJc�� :R�S���%_����>��^/��E���g�;a5���1%�u+�դ'.��A\g45����Ⴂ�3К����5�������(�`���#���YF��̄L��ڡ�{AE�K�pmbZ֣d�˃A�t_��OjQ��~��?j��v�"�,��M�[��so=JYz��<Y���C�i�����<\q�`��Ǔ&'���f!v}�
�Q������^��$�G��RF�l� �z�X?�@h{v��|�e�+����v��
[%�l��Y���h�in����z#��1�ft�%����]!�f95����@�NA<2�j�y�	�\\Ft8$���m� Afa���D�E�Z�(s /4��+{!��D�
�@��0:��{��$�Sa��A�Ц��[Xv)2u���~l1�OU!�7b~�?;�0��*[��{;��\�j���] q�S5�XT�[�N�@��`ʱ\����f#c+J�ֹȐ�ҩ�A|�ܓ���M�_�u�w=��ٗdx���orqϵZ����J��s����O���lm�<������1�.��¹^C�7t+��Q���R5'0��JK�zR^u��j���3�+�]�J�L�RV�v������-�tNcǶ�پV+��Y��T��B�� #���	\��3%�Tp����Lh�NN��{���ē�4g�e�:�4����/x�.�Ə�[NY��#Pbqm����[���}Tp�L��R�����$8������\p��kO12��u�V�!����/?잣���1A���}����AV��؊iǜ�H�l��y@l"�Ay���$B�!���/�7c�A�c�<; �e�,����_s^�ѝ���>�K����%LQAR���iuCFWx�
�=�=9�ྲྀ��JdP��Ǉe)�g?�1�Fٰ���?�e�XM�
��q�=���ڷ�B�+�`�����-�䘯(ϣ	a��/�Z��y�S�V.V�첆[ϞB�R(�h�\싰k�]I�;Ew�`�YEe1�Ԣ����{����Y[y�/�����aJ/�6��(hh�Y�*�챥�X	�\��������M���ɋ����`"Sb��x�"]dZ�� ��=��4N��S��Iݦ<��ؒ$�ÛcEk�#>%��9zR�F�jR�G�%�Y@�3�m����i��d��^��۬��,n�V���n�ӦI���2��N�dyS�}���{���u>�B��͞y0u�r5*�ۙ��˶
�m��x���/��J�E5G<��-J�����Ŝk���Ou��AM��t��Wk��i��Rdp���)��s�������6��+|u	~h�!f��c�/aC���
 )� �r��a��hL;�n������H���*4���v��n�P/(HN�;��[���hb���Dl�Q/C��0eZ��@�����]b����A���.���u|��+Z^>�wVe��.����?�����3�-�}B�4;@�f:n�1=Y^�x��(
�k�ڠ��#Q��
���z�&�7_8��^�/���|>M����2_z� Tw�r� ��B�Ȍe�u�A3�|�f��4$��d��Jm���f-=���y�#���)�{��t5f/^�=�����5��u�<�t_όT��sBq�;C�m4�6I��s���D�x1	p��"�9��am��|�?��m�I4�⸮���T�{�'��⹊�B��ol+~�S����H'�|��u��~^k[���ƴ.i9�����i�a����� Hkbjw?H�ī����'��*��HL%~,��B�LNHs6R�ce�ntM��[�h�jt�O�
$�L��!L4i�K�<%