XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����Ο�klU��:G��3�\X~G�W�R�SS�u���"\d���T�uSؖ��fv
Z�1��WΟ��T6�͊9���Ŀ-�5/c �3�9|��rm��g��ZF�Tl��َ'��G��r�m� ������i	|=2ol��v3G�c�Ĭ朝��"L�*j ��0ѥ)�g����z�,�&C+��5�Pz˖����������E�H��*&�:ź���������,ci�H��H�r���`琁!��Nӈ� �j�"B ;�Kye�gMb#�`BP#�߰�n:�<W̲�.$X�_��`UB���~���	�Z�y�V��.誘<��OJ ֝����C�iJ>-H�i?U�⻠5/a�V�"QI�l^���4����i�܏�@�rgS�[Mv�0�2� �9���Sl����g���b�Pm:ީ��V� ���3	����Z��Hq@ݒ!ڐ��x��ԛ�Z��)=��T���� +EE�I�
�@���iE���_I]��N2��f[C�6�=�S�I��������jȀ0Ąz�uj�m����h8	�)��F�(��:s�x��t'��8���i�%�tx��'�|���i����WxsD׷z\��˃�<�g�6�+j2�ـQ����3�ϼf1�p�T�#úpg��c^`�U�q��7�)�y��uӜ:�}�
��3����91�掫�t$��_���1�߳����݁'�ҧ��)��GwE�hyA�hZ-����,�/mXlxVHYEB    a037    1fe0�7�����ܙ`'À��
����R�&�1�<�]����
q/����5�/:_��P%���T��q��6_#�� �����K6o��T�#���n��&d�����F�}��-�5��?�nz8#�Zz\��v��F�֒@�0��ķ��L����0���|�[��}c�����G<���so�Q$�YZ�Q"_��\�D��}�䇈��yL���Pk�}��z�}[�!{>��em	�1��!��P.�}U��"�8Ѿ��P����}X-h]Ʌ,x������U ���(S���x��%~y�uPw��V���a ��z	�FU���zb����x3�������[��4���K�߇�-$eڇ�-{60�b��mǄ?T�]&.u5��1�s�Y�
�n�:�6�,
ibCx7JDH�}G�K�D�Qc�t���֒Nz���Ǐ)��S��A���↗rV_Xn�J3��֋yd�&4��TJ83�=\<��I
:�O�K�U�h@���s�������c��2���1:�XO^��۲�ob��ӽ�1� �!vr�g@�%RϝX�N*.�^��	E���'�~ey����m35{F�p��ZRK����f���D-h+�EU����d""gƈ	u�@xI\c��s{S}�
�=�wA�z;1����U�/��\��&bڇ
WFzFN@�`�~�ņ,�u`�*�q�x��(v/�^A��pJ*91�=�}��)[����EH�.k�ם^������"�I}��b�Ŏ,7�I@2-�
��p���.�F�I*��c UQ�Y�&&�9�'c����u�m�,���X�<܃�5��1* GO�)03p�l\DW�֠���V�a�E�)���y�b�k���
�q�g�nO��5���0��C���z�V�xQ���Gn�ڱQ�Gj�H�R�4I����5�� wj|�� y����Qa9{�`r�����!�
�j�Kk�H�b��W�4�-�!,T+��5��\f����i�A�ţ%������}!��ab�/@V�d����=ڟq8�RJ�0N%�@Ѹ�f�g"��3ߝm���j����UY�"/�ɥ�t���Ú�E3D����(C(�]����H����h�L"�_�=��0a�8���6b��8�i�PL�S;$���^�V�臜��)��dg�AZ�RsH�1
�w���E�\�M���Bϕ����m�5��Y�E���껬E��O<,M;bA�ls%P	hO﯀=Jz�؇F!��$������ֹ{L�x���^C������@K2����E��$��D���ӌ�Q���M Ԇ�珶��SE7�"�P��<��j0'��*mZ�(�)��P>%jחGR��z��^L5�"%�%].O˫N�4:��Jڄ�S�9
��/����i9���L�K/���nހ�������VE�p��W�ڑq��E�T�b
���ٴ��F��[���F��!&�5��n���f�%��c�qבCW�[�Q���Z�<Ov�mx����'I���Ꮣ�H�h�JK�?�~���:WG��ޥ���ͽqwP�OO~3|4>�����qȰ6��k(
1_�7a� ��,cY1�9ym��S��O����\�s�<���./�X,���7�E��P��[,1��Iv�Y��-J������ps� ��lD�c�rl?�:$��P��D J!ek�|��R�#�X�o�}��-a�V�A~_4�$�v���3WQR��bX��&�Z���w�8Q�,�1~�R�e{oF�����5����p�G��;c��FN�5���H�u�f������c�	N܂&��R`���t��^��r:<&�����צ?͛��4!�u�Z���:V�D���w�K��9A��ɪʰ�?B��Jy���J�����h1C�	:s�_§�=�7Q�7��]DR(���}
	L��-�1�jy��W�ӽ����Y�R��ʚ�UFB���7ܕJDM```dK�d�ю�oG2���:|�M��v�nByW�ZYت��[\�J�Y۝����G�]�!)�$_�֕'�#H���?�����=ųN^�91�%J׃'o�:���0=�UI��4]Hr��_J��i9�I`�b'�||����?���P� ����� ��	�ߨ�^q~����٭����R#���CJ}C}�z�ru-��kq�=S��:�h�bx��+��-�G�1Ss�џ>��*�i�8Z�a�EHѡ��yxI��0�X�{a���<�)��K�q������t�B�n��瘩�a����|����p��"G/E���o];���M3�E��bu3#�,�m�i�a�"T�v;,� ��#�&�6W��z	I����ʬ�:��n�1�R�R\{e���㗁�P�B�ehzk�M�pѪ������Y���y��JA|�pgL��1�-@�J���ȷ�c3��Quꃺr�����{��C�͏���4�.M��Q]�1V��>�oB���n�~خ��Ȯ`�]lQ�q�:2.@�-/�ڇ���$�����\�`�%L�}E�	َȰ�ֽ��u��2a��,1EU���zay x��i�����r�O���~��*Ҁ%�g.�Y[�}V��r�8W�Pd(�"}�_`��g������B� c�܃9"�զVd�);[�w:h��S���/'��ϗAw ��5�%ɻi�:�.�q%̨ �/o��1U������U�����Ӈ�c�=y6}�jz���C����Qt���K��1��m�0HtiF��ض�5���������/�����:��tG#x���w�9Y*�E;��JI���8��^X]��ҼF7�ԭ�*[��������GP�	΃'��qX�-[q�)e������z?⮅����%:��+��Z��R�o	h�� R��=d.N�7V���W�m�'�Pe��y��}TAcǮ_ŕ3��Q��}�$ޑ&.hk�kݝ�f�7t�_��G�f��hGO-�'z�x�;��}�p��`�S�2�%	o���37�9E ��c�g�[� _L�-4���
�Q^��A���Z��T��	���Bj�B�ز�ҧL���n�v�W��s@.�+i�eB��Ln9}��=h7tQʾ[߷rր�_��/�Xu��T=-?����(��Jz6��
�P l������4��)���e���J4�7�.�h�!��S���f���fwьj�b��qTap<.�
��ג}��I�s�	Uz�w9[<A���٫[��@S�:ԯ��b+��ǐ�Ob󁳼�%�EqA�G�ʀvOD�)�_�aQ=��yN�?^�'���ϼ#ͳcI��9��ی�@�"p4*��<e��-3�L�]	�<W����5W�� Ko�ml�8�8�y�˻ŉ#�� �
�����)vdA!e�W:�z]Sub���2�'� GBj�27<�8�`i�޼͜�B!�\-䬄C��P�Μ0�K9��(Ϲn��k���Ȧ��,�K-�R;MŢqQ��{0��~n��RN��}��f���^�Ý�㛚��7J���+�����u ���a�����'b+}��D.��.�c��I�����>a(s����j��ĦY�ut�?U������:�Xm�X=������o�8)�"�2~S�g��3��僛�[l������������<���;����hy�rੀ�]b�Mz0���
�ū��X����n�V�� =�ed�_��sʍ�m���d�li��}���l�|5�Y�x/_�-�Ɛԍ���)+=�S�ȿq��W���������>-%ΒG5�~�]��8(����n���<{������08
r}����]~�����/�-��D�V!H�O(����x�b��xX�7Y���W4���#RZX�ihy�����j���x�[I���`3t��{ėG9�p��}��j�o����)��g�JtfaPLh�Ѿ�Hso���H��U�v��f�d?����gr��V_�8
�Z����d9��
W�hZ�p��$WuЏh�2�3� "`�����,�����2�F.���kD� I$0P�d�)/A�m�(��<��D�\�R�nT�ؗ�-{���l �R�2�������^3��,%f�����]�j�	|}��n����b��{��$_7埱��]yج[����n�K���N�R�ӻ���tZ���	��J�~�{�y����sr�`J�c��x>O��i�}Xl���z������'��(�wH�˞d|Wm#?!$ߞ�ff(D.'��O7�F����k����.:���1��mD�G�������,�I��W	9Hp�w^���4l�v��g��j�I��z�-�:�|d�k���g�8�&�;Fs`��ĭ)M��1ʡ
`�#H�T�N��yߥgaUY>D�&��>�p����«�e~��(jdB��y\�0���]}}��)I9�<�Hʌq���xQj,���.�9��yCe��<$[�X�*w��v/��54����蕯�Gb?���;3�>W.�L�8�2};i ;�ॎQ%�1�.����=�c�B�{Pq<�X���9�����z��.�3Te���[+�C��kR<��z.`�{Bˋ�8�������Z^�Ћl�F��C�S� �q�k�S�8'$�O(^lꧥl?��H0�ue%ć'���K�:�T�Q�&z��q�R�<*%������6��li�P��l�j:UQc{�Z���h����-�ŵ8�%���<!���֕.�8m#	4��b�A�IM:[S9��&<�4��-ӟ� r�Aռn7��Xڳ%Naj�B�2��s�9��0���H��e�6uW�9��s;������6�u?N�}�O�{�&�;!VTI�[H_�r�oH�B��O�C�d�;�@�Xzb?�\�h���'��?
����^cS�MFn�my���j�1u�.�����Ԯ�����IDy��a�ז�.g��S�N�q��-�֕>����ZA��{xu�P����ĕ�G�OkX��*)��-3i���ݖ5�p�c��$Wc|y�W��f89r�7��tu)^I��[�̭`�����S����[�%�>�8�v_��p3 �f�#�֩9*�-�0V�7�&8�؂���4�x+���3QF���B�l�l(	��v8�jW���
J�M�;��S�/<}���!yJz�
jD
�-�.z�?� ;7¢JB�����Qߨ�r�zY���0'��Ho�$\'�-iJ;  �}1��F2O���#ad!`Ϫ��bO�:������U���Xw�?ӁO8�g��������T�Z~�<u���^y�oE0m���xF�L��1��Q��{���'�M�y\8����Ť�rdպ�E�����q��N[�Q��hO�<������,<�`��x���.5M{�i��&1��d�01�B2��=�T�~&KGf��keLگA �����U���Իp��m�?�N�#�C�hՉƗ���}mlO �������^��1�W}�y��FM��)�䏗\�MVRw�龣�Њ���Q��[Q��v��RhY�z� \g���T�1g���7�(J�S�Rߓ����熈�(�D�n���W���W�V�1��U��iC��Ⓡ�>��e�8��s�Lg&��*�X��=�$GU��ϊ,���@�?o�����&?�A��$����;�?O�l�`�Gg�RX��+/��)�=�8����x�O��P)ǚ��ZO�����R��R ��/�����G�۶�MjNݥ�Ep�'y��+g��R�8���4%B�%=�����y�`;d{�Val�>6s���n���(	�;�f�Q���/z&4
~��꿮�.c��M��&�h�Gۭ<"�提�Afz	�h@�Sy�2��Z�'�����q��q����XV=�O�]�Fj���OAf�>�n����5���b�\�0(^u����9�U��v��*e(T�Pz��N��9��J��㞚ͅu6e����ee���h�4��1��2 ���(��}Q`�ǧ��xr{D�x��e��K�'E3>7:'Ë�a�r�0����"jE�:WΏ���XF͋&�L��������2Q���ݢb��(�*:��т:U~Ez�a2��`�WA�!<s"����V��U2���������*�����F��fkv�\�����$K�秤-ݽ/��P�+(�S9k��%{���������|'I�o�QI۶)3%X�wֳ���wn��~'�d�<IP�ۋ
l���a`�K2�]�[hn~Aj��e����O+�p/HDl��#7Z�-����)�v\Mu����O�΅�%Y6�4��v�����m@	�V�Yb]+��]�ˠx��<Mp���L���o�i	�B}�`�vG���1J>�G�1+H	�nN���wtC`J�6\	h��mˢ�����t��֛�#j!3�k�q �'Gh<���!e�>�=��U-F��dW�k¨�bݛ��A`����£����X�{�)#
>�����:D�4�|��N�NI��x/�M�BX�Fd��qw,��|������ZMh��W]�(�V ��J� �R����`r�Ӆ��سn�~�.�`X& $_�'^�8���ߒm�j�x.y���-,׏)��
�R���Tx�I@���/��x�#�k�),*G��+�E�Ⱦϯ<pm�SM?�"��h4%�x��l��=��|I�_��"�\#wF��s�aeڵ�Y�R�N:����_�!�# ����=�h�ۇ���'oqT(s5�J����ȇ1����h��Dm��u�Б��`g,� ^F�ꖈ�Ԝ���>�.�򜟵����J �����ѵݸ
��<���t�P�.6城�`RY��0�p��Z�S�a1�	;�~��@��4�����#�co|"��Ɲˁw�Jx�Ё&'i@�_�0+��?g�dEn��Q��7v�r���
EOn?��ٷp�3�jDai|d����r�۠�Y��ߞ�,�3M�>W���)�T6���3 AH�^P���*W� ������W��rD���,�v������q�Ȣ�ͷ1�7��/�C��B� -�'���e���PywN
��;�P����1 �'���A�оZ4K��nj�عQ��Qv���.U�� �'�,8�Mz�PޣB�����P��TJ�k���ݽ5��tY�I��'J��1v`_��&5h[k}W�	;�*��r�#�v�pH��56��+�C/Mx���y�U�EڪQ������P��*Ȝ�$�e8kQhb<z:�����9�#}�N�g�[Qc�e8��Cc�`S�B?K�x�ل��|CN��QPUJh^A�-8�~�I��|��V}�G��;�*�,��pL7I�.E�q�?�!oH��6�{W��\�ij����ǡ0NmW9��q=�߇���$��m,��ג��Edai��%��;C�!�� .�9a�[,��hV�6 ��T�:�zNdgo�7�7UҤ��3������Ή;1�8�(�*�hE�K+�X���ۡ���SV�.^��))>������뫛�+c��XsLUw�%ʗ���{z\Us�|���H|�~�d��.c+ϑ����۳��UR����{8�����O� ��K��<b'�X�[ߎ�
�?�QD��A���p{��۱��p�yBT Tӓ���@-D��ByN�`ӊ9�A��e<�(X
Q��3_��Q�@��Z����� ���\Vx����s7�<�s<sí!�b7���?c�$�5v�"��p�`�#d���N�P �a�z��[ ɦ��j~fh�uC��[���f��\_�Y���mn;[�P��ܐ]�`�I�EGXz� %���U���n��0W����q�0�i*������瓘���1V]�nU�J�YEE�~�`�+}g'���a$�50�s���W'�9"ҩ|�B�c�TQD�/��(����X	�)�P<��/I�$�u�!���@�xX�\�N��1Qk�6�Z�%��%��c�d~$