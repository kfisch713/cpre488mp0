XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��iq��6UL��Cl^)\�p=�� �����)��0E�����]M��p �n���Å�,��$l\M�C�"�]gw鳊�#qL������?�ֺ�vQ6���r�ʥ8l��ğm��n�H��'�M9V���F�|R�F���xm��}u�#�f��k&��R��I��������V����"1j��<�E�JAu�'�X��ë����r�(c�f�-�?�(��26�U�[�d�q��8quȯz/k��ن+FI�x��͸�X��$#)}�ǥʿ�d�B��Q�E�i��בC�ky�7+���i�����X<�q��I�B�!e9�D�{�~�g}���^ܘ6)rx\��y������%ķlf m�HI���xw��_g�7�����L��w�e�N(=���L[��˅��O�ۻ�&�K��9>�^B�6aF���g��@y {K��`x��3�`�*+*��K��C��F� ��!��'_����r�r�����P�'��&.����a�5��&�?���{�*Zb��O ����G!Ү�g��^	:b�5��.�����,��ͬ@�XX�@�nI'�z�o��6��z+��:�8h&#��=�@�X|�ތyO���N�a�^�r��w����,��|~�[?wa���;�< Cv�s�o����fDig��K20L�;�/�*�%�{��`:�^�y���X�������󦼲�cC��L��a� n�s�s�K�N�	H���'�k4��n�nW,�XXlxVHYEB    b3c6    25b0JB��-�Պp�U�I� pr�S�_#��ޯ.9�&�0@[�`����������\��1�(Rc�q�e��|+���;]x)�	� �,��\T /
��ɗ�� �Y9�䆿�Oj���V������n���ɯ�dW6(_Pt�X�ҮS��o8!Q��*E�s9�)$�;�����?jr�e�z��Q�ES,��ԩH}�@S��o��G>j�I:�Δ��Q�P��V~�H�jPH�z�y�d8	�}��K�K��a�$j������)	t����<u��؜��	 ���f>���Z~� ֐��������#�'Nt��o<DR��Z��Py�^�sA
��/�0�{U��Nm�$v���]�5��ʍy�G��DJ�)�ݾW^�@}�V1����jK���1S�(�b�u��7�v׋�����=��h���D���z�GX�T���ŢJ�;-6��rl�(�0JI����Q�2.�<��iC�!���8\�I/ ė���5�B�sx+�	I5e�}(�x���Hx啧{��
�� 1�
{�[͠d�5M$�[��_eu�/g[�[ĐwG�G?',{;���aU���yc�/�|=���t�+���o!Y���=L:d�*�"�zWdH�]�!��Ur�ڹ��5��I|IՑ�f�2ߧ4��2�������}D!0�V��_����SKQCi���e��p/s���H�����תS[䃈�]э~r�!_���[=��E]KIXlmʈ*>0�1[X���H^G�"��x_����cG���g�#�&����i:X��$��W}3��v����'9�ai��F���� ��X�0���Lׂ�"� !��i�����s����" b���Y������-ݼAO����^~v�A�.��-^��>(�%�y�a���|��fD���+�"��	ۭ�%�{�pH���o@��pB��щ���o��_#�tA��)��t�+J_�ﮈ����z��5YI��U�$/�@>4a�Z Ȃ4��.E��ئ��=uj����g�޲ȵ�{�� R�~�b3�4�+��-�|륿#�"����vU�Wk��G�[�vA4�+mW~5��U�<�b��右�h0�K����?�.W-q�ckk����jנT��u�ilP\�3z�+�I�X�>�N)������2���o��q�Q(k�Q�zġ��Xl5JJԦ�.ql3�=��A] �6E�3��7�sɬ�@Ӹ"w��e��������!0I��P$׭L���7�
❖�;����*_�&�H�O3����j�{�=��' ��=��-ek����S�vڌ̐.��E�a)S|�z(K�� ��J�忮 ��'���?�s8/Q�3�.^����O�oD��I�Jc��P�?̝��c搊P�;�DN��3ߡE��otg{Qo�8� 7�T��h<��9D#�����������%��UG�ߟ��2[䳛F��5[�>�6�璙[���z�� �J����yd�w'm­o�u�rZ1l_����e����o��M�e#�!��¼�7�R�����Uн~�~�֗��x�D�jw����H�lh����v�by�	�����[��h|��ē[D�)!��IP��\8�3��8s{��� 
�*h�W�������/��[�{H�ͣ<����3k����鎔��{5���&P.�R�49n$��DwrV>���_	��m���S7�.�
v/ɇI�tb��Q]�hE�C\���c���6X�]��g2[L!������]�%�J��~Ym��.�zJq��n�*a;&7�.ۉOQZb.w,)f�4qݵ_�Ϋ�5g�Ï�ial����ř���P-��l5��8`���9��lXR�W$֛��M�ȉyR<��'r4�#,u��P2�'����"��o=�ъ�M}%9��;.��I��<�P,dWnsR��p�*A��kH�����5W@%z�C(��{�5Yx�0#xxO�'�]�3�Q<���J��-����F([�ei[�	���Olg�\�;b�ΨI��팅���aĩ_P�h�HMu+6�9s�BS���χX�+���FVE������ ��\��<�1�7|�
�����:(��-���K��v13��e�퇾�$��F1R�zq?�p�m�+������Y����ײ�ҦdG�(��l��k�����$<���-¼��	mg�&�ͪu�y�C���C��m��@ـ�5���m��q:.����h�'��������h��h�WZ�B��®_��J����xE򋶙�P� 8��^2��_�'^� ?=�Q��Y\��ˍ؎�����J�জ�p���b��G��M�昮�.�����u��������q���=��V��JXrԤT����`f|8Z�W.�l�wY\���Y����#ښ7ge�*۽����J�^۽b�i ��\����)\�@�Ś�L?��UIC���[�A�J�"�v�c,�ϒ�vR�ދ�v����ey�x<�a���;����y(eL����.t��HH>��fޖY����b�+�	C�A��c]�eD�*�����y�®�#ؖ���nf6¸��/Ng��Z��e�.Zݑ%b�Җ洋�@P�Nf�����sAן}���\/�L��-ηc�"(����,���?��S����_��c?�G[���f����&�������Ν~5���#P��i�MU��c��%	}p#Ve(�[Ϊ엝ɝt&g��22#�{8��+�����;��b.���6��x_vI-6]K���&�K�:�t��[#�@u�_}ʔYo4�X���^צ������w�����tv�ַ��)���V|�&A�s�_Ǝ;[��[�����a��<	:�'����o�50o?!�tz��Z�i;vtL�R/�V:���D\(���W��3� y"Ҷ�[�h}�UOl|Yr���bZ�x�$���,6v�u'ΥC�hX��%_� ��c�?�	��7�^�2����0��8F�"w+����@���
V\e~v�Y�]�ej>a�W��`�� �Pp��I���W����4�6Ԣ+��vLB��DĒ�UV�o�t�H!�AFC,�V�gzY�U2��?Tda��JUʜ�(��
c��@����bZ��A��:����'b�~L6o���C@���b�H�J�Y���"�T�����	����ea��_*H�pe�z� ��{�i�8mQ�q�/��q�boڣGSק�������U#7d=��qᑻ���s�Ir�������,�n�PW��J`�=�q��k8o	J���zT����u�V�(�3�~�a��2�H�=�DVb�_K{�M�Ӽ��s�栌�n�Ha��� ��e1�ݪr�����/���������ndA�Y:��\b�T�\�� =�u�)�%2�� W��ii*�L���v|?���.v`[epZz|Q�{��������//.���!�k��k˗�G���[��\��>I-�m%��<TJ�H�����*�& ��ZS�"q�S��kj��T�d�̍Kl�t�D�`�w*��?�:���������Wㅩ�>�g�����@�o���!V��Av�â��e8c9������`sZgXKb�A��;�OQ�AfV#і�dN �0 Q���6V�l�)��k@�LVO�"��w����^��m$���z��Mg��|� ����l�'��P�6�A�����ܯƢr�݀P2�{�0�np5<��i̔D����=睫�� ��'�{�-��n��9\�ͽןD�����S�&4�����+����o��#�1I��e`@�i���|SSl���Q��7pd�?w\X�zl��UŃ�U�*ƶ���`��.*g5~"-{B,薇�TT��2��c����8L��Q��p��ކ>��|C�O@"���P/rQ��hw�FB���QF�n8�3���r4Tݾ����M4�Xd`�#�_`��7�zE��pO���hGr��`�@��hen���W���� q���S� ��-PPn��߅��aH�)���F@D����zw����>�M���~\K�FD�m�C՗Z'ih��ڙ���6n��]�F�K�e���b!�Ð챖Ꮢ�R	��ޠH�`�Ԏ��"�tFD;�Cx2���)�����׷~�^��
��-�O�DaB��(�����S��r�2Ԗ��|�w�ml��3��܄fo`V{ :1"�5a�I.�2���I-�Pъ�'�������W�v�����H����JU�hN��C�Td���.���a����A�9jw Ԩj"2��:}5�k~%@d��yXq�W�p�x2���a�(o� �x%��: ~|��Ŭ�����S;nW�� b@�	�~?.:��u.�)��;W6	э�Ylo�����A���sA&[*2�=�'��r��x͉-�3\�Js�ѯ�!l�������6�X�I�&]���C\7j�n�ʅ��T�~w�{��&X�G �V��%�Q�0Xv��	t|,��F��4Y�q>�\_؅�`ᚇ�aqd�^c�t�����-����o=�;�v53:W�7��Q���'�<�y'�2���O��>l~�v6:��,���AY��	#�^��Q\���c�ß+��ƌ�-6���i�A��h͵�<L���a3�"��*�v��N֕(ek�G����L�ܕ�$�M���6�"C����� [Q���&<�	���sX�F�J�i1�]=���m��JaB�{�d�Tյ�(�,��k?�R:.m�i�����Rj��L_8�&�,�EDd�S<��vϺ��}y�0��z���4�!�%� _d�Q�/�/-�q0����z�w���BK���&��}�褰(Uo��kL�?ە}�6y�sx��$��ᩱ����+���Y�8쳮�\�=f��O6�����*����O��In� �X�	y��y��h�̌F�9�~������d�h�Iu�	E�P���5�!�\����7�r��VC�]hK4E��>��A>��J�ǋ�&�ӟ�\:�E�F��&��&c�8u����!" ��T��Ay�;[�saS���8��9+����Ċ�Ȕ2�s�5��2��G�M����ͥ-�ǉ��Bq���}J'�oG�;�)c�.�N�%��Ą<�"苁�JG�D����gQ��7����m�������L$�%�w����9d��M��꠶5�̑�O'"D��]�w?�y�9��$�L�d�;�|��ȺUu����{�5��^	��"fWm-�.e�52�7"�G5�0��Z�B�>f�?2�҅>�y� P+Ĕ������c���d�X�B�x�\`�������eW%υ/�5i(�y�������ֈ�B�A�:�ޞ9u���W58�%+�Nz5ŉ=%�d�`a��ؐ}��{�s /��N"��y�c�eҤ���@\B-�FF3� ��?x��CT	A�ӓ R��<~�w��9YGtG�x��	o��J�$�M�츊˾����#��\k�@��]���yT���B��[����eN��8}O��;+R/��`�,6��Ӯ8ZaZ�%N
��rM��-'�`�"PR�ts�A���+�j��k�ˏ�:ܣ�lť��Y&�*%�@�|=H9�ٴ��Kt���9�PX]@;+v	4��@4��q� ji��1���t5����,�>Ǯ�y�a��U*:� ���F���훁SX��qJ����4,�X@Ϫ�C��?��v�&�yVÏ1�U"��]ރ�D4c�������ņ�]%���9TE���\�L���o��K,~��w_#�5b�i�rS�l���H�ߣ~1u
�<`���'�U�ޗ����L`2�N��O�Ꜷ���5��\�*��+�>�Ab(Aǘ�����q���,�h��?Æ����������`���,d�ቅ^��)�(���oc�ɓ��=���"(��i�]M�E$���Jo�7�E����� 1�y���b���<x��ARq�d�I JZ��8�@��B�7+�z蓑LC���>�ۍA����˯���ul���ˆ�G����BhÄ���n3Ȃ��H,�� ���1v�� ���F�]�'�
�oa�����dƆ���|@�$����cl��s��գ�3T�"g��lո�P �(�և���[I)6�����K�xB
���;���0^�M�� ���2Um���W����&�\6��ݐ�v�� гl9b�|g{���:<�X%Ļ��h�B&=k���_�B�S��ٟ������փ��g�5a���.�����Th��@
�cY��C�kD�k�h�������N�D��m0��K�����r>/�oy��m�x}Ņ� |���@�'�\��*CIH("�^�m5Oʛ��lJ�x��� ��'@=�f�((F*H��֊��p� 8��+��D�$��b��w3�9�p�v<�3](n�P��b!����Q��=�"o�����!����m�cTu:���L��+Ώ�n�XZ���<��D�d��1�-��c�Y������fޟ��AYT#l�}uP���݉�*�
��c޾��,�Q����)��tU�UȐ���ȏ�a7���| ca�wײ�`6�F�:��sݨ"l,�Q��?D����N1��o&$�+��˙W�3v]F���U�*G7<�����Sxу�PU���
�����p�񵮵EbzV��%1�}���Z����^Y�S��ӻ��W�/�^����Wb�Y��"�$�K�JH���T^����E�\��������R�*!�qנ<6C��T����5xgܬ06�����]-ȅ����#�[��r_��.b�
���BJ����65�<N��Yk�gB��|A���Y-��I�d�'���$�@�2%bbpݏM1�hPA�]iP��^����;X�~J+O�i�G�ۑ�7�����s��z?�",����;�a�?]�Y6ʴ~̽�}5�n̲��v��Ҁ��Q�[��f8������2@����k2���}�|�d6"Tg7��j9�^þ��]����^n�)��y���F��9�yXk�*�'�Y�g��!�=�vYi���Uw����*���r�(S��R�XU�G0��q�����"�L�a��'�	\n���z�������7Bc���) �9_�f6�Y���>'��{J&-�:�����|���L��ˋE�N�2ń�p^I�L��x	y�[ݸR���N�/O��"�O�|�
�*�r*,'��1|&�h�����sy��r�j�̅@�h�/�<�d �A��:y19�	PJX^�|��R9�w,���:�d �5o&�� �<鄑mX�������_[s�6ş�"�X'4Tj� i'�/6F�z�I�ؑ��x�V԰,=��h0Cj�����������%����	�ou+�MX���Vx��g'�Oa��'�2�-�!�ɭZ��w��ΆȒq�(�ɓs=Kbެ�6L��Q�2e����J�$W�Qb�=ڦ���L��hN����$?��>2��Єp�k!�D���~�k�[�s�2�R8�����'';��!A�f|����tN��k.#p9�����8E��D���Y(�A�W.Aߘ�x�=@�##@D�U�֎��*�l��y5D$�� �1���(��?��d�2��������"�;`v�dLeOC�]V����q�z�hGN�0�.�T��af�>���UDe9[2fг������Zq~�x�mY,N�bP�L���3aIһ'N?�I۝E�j�(����b��#(����,��S�ȧÝ�)�[5�8��/ F^����0Y7vi룃GV<l%ߩխ�4�[x�᳜���NS�������Y���ޤ"
�|h}��ɬ(�LZScՃ����r��铒�zѤ�xY��Q�Ә������:�F9m�pD�����=�sDx�Іy1X}�C��G?Ɍ�g���.p�a��s)N[J��c�2,�̰.l�渔W��K5r���<��V��2�~��&��C��|��tB㐩~4Q���*P�U �-� �g�_YG�^_�vlʊ�o��6y����s��Y�ߝ�
!���#Oj��+�{S,ސ4�kw�� E�wT����cM�_%�G�~� ������֊J�8ְZ� �By@8���F8V18���=��H�=���^�Z�p]�by:^ ��L��(5��[�y+m��������K�K:;��|8_��PG�dH�K��:���C��%?��d�$.�������.$KX�f<��9��=��p�s,�.�_Њ��a_P��^���ty@JڲD���s�{ZX�2oZ�"��]�(�kl��:�^� ��/�5�t�BЎ<}����L�EÑT�'��B>�Y|�}��$�n~H�_��r��;�V���gzLEE�]��lɫ
 ̢bWc�~hq"}��YE�io�tۀr�N�k�-����D\M^�i��Ն��GSnL�Ip��R1!�L����L��l��e[U?K]��^%}�V�m&�0���/��:꺽��^�c<�假�4wF�qF��Ϝ�~���n�>W�F��c-��G@r��f�uIq���ȃW�>F+�N���:���B���2�ߎ�1��Ff�(�C��X	��K;�L�ULÅ�G��@�5-�W���Vq�7"�!]4��O@��5��#�B���ȴ����.ӊ���P����TN�k6���c֣H�HGr��񛸺�{�p�V�c����oU���mK�����%���|��eN���-ɡ�QD9�[��(B�/���1p�S�E�S��*���kxA���Oz����������+5x��[��(أ�����i�s���\���J#G�]X���W $k�\�%�yrښܴ���Ž��(�D��I2�~�΀6JFޑ��˞w�L�LR÷Xa��!ٺ�D%
���Z�O8&�M��Xp����&��P�_^�.���?��Z��
��׈X �5/��TV�����0i��4���Ҹ�_� Կ0EUJ梭Dk%J��Ǵ� QG��GN=�~�tJ�|��X����>��G�܀B��6���"�u"�2��`ɆU�̍ ��$�ZV�ē��J�}#.�}�|���5ÏL����8g�B=�"�F���vE]!q�D'��u��kE���@NmJ;�~�xci��J��y��1)����tґB�|���	���c��\���iJ&5�a@�D	 ���zA܍%+~^�@� �������`5DJ��FXM�6(cW��`G�����:�,.@���X�R�̘!%��?��*�3�݋j��s��}Z��\��C���h
L�t�TM����P�)���qH@�qS�GtK��1��>0���$0Q�kFa^�Ҍ�]�"=�E���L��Wi�LU\����3쬻,�$�#���e6=�H�Ե��GeZ\):�Fk�˱��"Ⱦ�W��y'=���.	䉭��g7���l�n���^W1=g���j�[�o�D���