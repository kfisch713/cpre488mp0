XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����3w1���E��It��E	�B��v]����L��<V����2�4b�5��}G��d��?xy�dн|���>l�Ѭ���+�JH�]�a?�COj��2�S������=��8�&){����ä��[�[ϻ�`
q
��cYjc������j6�6;`_Mo�D�%�jxe�H�S��	���XwJ��k�����6����8>n�E��B���i�����d����4;�郈]�!~l�K�k��M������mZ�n��r����KR+��_�oNP�w��eXd��e��8�7:K�L��:�k�U��9+K-<��4��ܰx�.��e�M�'�R[K_hf��7��'��L�h!���2��[�����ꊀ�y:ڛ���5Ś�"��W�B�<m������`.3%#@c��ߙ�L��1j�/�k���[+w�@P-vUbg�����떻&&�ϔ��a���k%�Rڗ��;J(N@|��ԝ�
�Ca+|�:M$�h�-;�8C�H��*���sm$����v#����K��GL�gO�kj-g����EQ�Iͳ�!-�v����V�~�iSY�T����}�R�|����aGo�� ��G|����+��9��5Րi�θ�"«7�2Iߵ��ѻԥ뚕�pL3:I��j�TPP�!���F��r��k �h�M�/�l��7Ee��ߩ��`�^\)����2O���F׻�A1b�� !鶮�\�
s���K����t�ظ2XlxVHYEB     f6d     6f0�"`�����b���x�ja����m|�R7`���V�V��G΢��*���Ʊ���8���-���W"4�M��>�D(V&��a���^�>_�:�v#�!�v�$D����G�7�w��ۉ���)��H��o*F����k��j���N�(Ⱥ�f�ځJa���f�h?($#ބLlK���I�h�5^?���-Q?4��k�%��6t��i�p����g����Ԣ��}�0Q�2
/!(��OYh�p!�{�|�tEgL���g9d��r�{&e�"�\7��˼r@�H�j��d�1a<�`K:l�+Y��6��L��H��|��[wx(\*�bN�	�7�c�~t Τ���BetT�r�ٞK���yLҝã�g�|0�,�E�fc��%s.}w��냲V�]�[ϡ>Ͱ���(9!8�)b l���&Vj|�VS�@`�kICN�l՜1��[�����I��5R��%��}#���xz�)�SR��V�N<j4�-�qԻ��Pw�y+�� 5�'��P_�Ty��Md��н�d!�OUc����Q?ЪU�sY�����n�B�O3K�!������_�G��4`y(͒l!�,��A�CG�2�_3���;�f�Ŋ���M]��
]��ʈ�(�@G��S8Պ��죀��XU��Z�w ��`��*0ީA��)�m��<�ސE2&�	N�9aaS!������+Xܙ~���l�`�L�.�Eˢ�[Ż��>"�@D�n�|���-I�����9;j���������3�!���F-ɍ�u[v]���Ѯ�rdx�Hq��xP+��,Jo������Y+c~4|a�I2��q�MbF�&-�.//��x`�,9�[1 �����u�`Y`�N��r�2K �{�$d(<9I����J-F$a�Bo2_p���@3��²�[�j6�_���O���k��ij��70s�x����b�G��Y}�o8�����:C�!xZ�yE�!�H�3x�N�:u9o���zZ��
��gf.R;�
XU "�v��f4�t$W��;a�ȡ�`f��ez �~��������4������������>��12�ʾ�^:U��E9�>U $NI���ȵ-�~|Ab�B�C�8c����tK��M����1�X��!Cq��������/��,�[�yɨ�p�uI���x`fd#�a��n؈;�S���P"�?'qE:�����7�F�$��5�u�a8�]��li�Mn[�'��z��2v?��V;��i�C]��@5GK<g���C����>>�"���R,uq�%v���ҍ���m��T=�&���N/��������A���������9:(��ϋ�`���u�X��s�翬�Z�{��O2\K�%�)r7�(p�;$@��q�?=4!�1X��4�#��O��5=���'��kV �Ip�9����9�ս�v˯���S�-f�Ɛ�S���NW�ٸ�;���c�O��Re��
>.|8�溠|��h�"�f�RW�*w�j��-<U��l���5�|�F���r�0��O&��k���{6�#�rfQ����r2��rż���J�!�Q5��1�}�ǥ��zD@������sB1��^�3���p��]μ��\��k���Pt�;o��f��~X2/5 �"�A���@`�����(�ۛ\��Či��7���hG^Oxp��,�����,Ϫ	G(Q;`Jz#�i�ͮ����#�H��lT�vW<