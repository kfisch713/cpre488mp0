XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���KP8�pj����oH]���]�>D�lԘ��7�;��
�I�;Q�{�W4Jr��=��L�9ӸP��_{c=�pg%t_)"���F�D�Rp�i8!u�p�����Q;��'�:S EY�������K8\z��|�|���s��P�ز���6WX��L��y|��?�fH��mL���(V�M�v��A�|ڢ�Lr(Y~��j2���gB�e*�`�� ,sz�2~����w�����,;�ڄ"�,Y��V{��'��柏vY̈́|�H�&�����W��\A��>�0
V2��0]+��k��ͺ�������A3���%K�9�1�Z���}��m�fS�mK{�7o�mM��jM��+���<G�X���x�{C�����8(^��V���]/K�|0(6P��t���\�Uj��N�������Xp�E�GH9�޿MlG��l��0�q��Ey5u����e6��R#q��C��p!�b���5�M��:�֟�D�nb`��u+b?m8�yR�G���+l{&gj����p؂�U#�̾	�O�=��٨�_��d��uEs|�O\�IѮ������a �w��X��<���/�CAJ#m>ݿ�uaol|�Qح�EL~�)��3�9�n�U��=Ғc����W!7�������g�Т��R�3����ͳbi�M� ���jxI�-6�0�J�>���3�>���Y�%��l�XEF�r,a��;@��Q�b�C����uȖTG��|<�����'�XlxVHYEB    b3c6    25b0QZ~wq$�}	�@��̞(����&����*U�W㏶��>W�jidQg�N�?_�U!gjL}y2<9we�.��P�/�L;��zd�$2�B3�&<�_ ɚ�j����a:�s�%'��6�Up�=V����%���-ҿpB�Ȉn(�'P��rY�V�uk��ϕ�j"�J��4�mn��]�����(���Z�8R���`Ĵw���o<�k{UN�4Q}�k��c��Qa����r�8��
/C�lߙ�P��zn�4�Y�X���7Y��ӐR	4%�ڒo���oo��ܯ!�f���5I�;S�K�&EΚ� ��}
J	*�c����H���P�.�s��g�g!F �Q;ݭ�h�(3��Qj!F�[q����w\��r]h��r%��n�������
#���=�}��Ħ){�B�X�D$Ii��{�jW �:[�-H��+(Q.U����Y��ovС�y�i���z�䢡�e# �-ֲ�
���.J�F�?�j,g=��ޡR�y�ͬ�{��3�{�F#��&m_�@<�ڀ� ��m�6Qm}�}�4���R\=��uU2<e5�pe����{�u�P7]y� ��c��4{Z����z{9�u�ZP8ਓ6�Y��]�R=+^�VʼR��<!��r����xw����oVs�٦-p����\nd�-��{1��/t.�_F#��D?�]_�Ce�|Բ\���N2�	�t-H�X���>47��-�zK�u p�o�B�TW��N$�k��+�<�f��%�a����-2�;�0�2�u�����bw�y���&Pf�D�����Uau�<��;o��f*ѹB���?�8<3�r�c�=�.��k�g��-
9�9h��bG��?���ȈK�*�����*7��kX�W!�^9q��@+]A�zF��:�����������/��`Ӝ�T�����DH�
�ю x�͂��L�
���ٺ��p۟q��Ŏ���Z�����D��s�6tFp���Y����_���_�hTwm�Wcr��0~.'u��,�H�s;����a2E�QKSѹ�'�ͥ�?���[�Բ�\qþ�B�ߔ��c�9e������Eާ�U*��d=����e�p�Xx2�0��TB���Ƃ<jƹ�XI	�۩j߉+�ʂ 'љd��t�����9��_��^���U�p7�d�"�
���h%5Rv��5f���Y������D��&Ә�S�N'��j��:r鈋k��.y�7��{�]xg�U[�+�~�
U)8�K��F	���Q�$���"!���t�A�<6R�+jSu� uP�H�Ս�����P�u4�O\����1����F�vC*z�9K�y�5�S�rQ���w*2&M�0Ѱ^�A�<SGݖ�`�R>"͛~����m�oԛ89�Lii<x7B��*��S��$U��~5ddB���*XC�d���_��=Ҽ'��_?
J���
��	bih��o�H/5$SF3荌z�q��Ա�:�����b$��6��g�/�:��\�u[�6�k�����R%�?g�!�A�����됔����'[mၩ1ͯs�Q�@�{+9�� �W���&";m�Z�A���f@�*Ae̷��5����K�l�X��&RC4@�Ȓ�����E��/��[���F0�9�]����'?�
b�!��u؞��pB-t�@�o���7K
���y���M���&��{��D�&�*����rp�sr�3_�&k �w�5n JF^AG��9)�`Q��,�CI_̈́Dc���:n{!���o|ؿ�o�[�j8n� �����ׅ���,-�9'���;*!�c9�G�a�h�5ʊu+B9-<1�:�|����s	�@rX��t�{� �V��Q�ng#'؝9�����V�8�D 8xGA�F����;U�f^[7"_k��9��MS�BF�*��_�LЇr�Ys��h�$��!>c.�xƬ"�#��8�>��`���c���EC������������cSW�   ǈ�p��*Ę\&�0�\1O��ds+�'��7O��èr:�Uśy��"�C�ڂ|��1���3�G2�%����~�?�Q� �v���D�fu�3�,6����_n�%|�Q��Qi��N�^��S�'����	m�'��L!w��Kk&�a�~�T`Gc9�	ɘ}���h��� �r�$_��P|!0�M����M�UFb�)=ou;����(��U�=�0p�I�����+�<6��T��j���_:q���ʌdn�k*�ä���w���A�	6+P���FX+��Wfϊ�
��!�xxϵ�ljK�p-��hT��r�|HV��! �}���S���݂#���؏e�zM�Ƚ�,Mw�=�Β�W���>QWAI~j����7KM��I*��L������#j��V"������ќ���%���S��
Y��ҤƎQ����մ�/���f"�{?z'jhBK}A
�6��� 0I��bd�Ic1��~��5��Z�"��ë��*��I��r����{3f���U��ew��������%�XN�2�Q89���W~a+�P�E����v�L�x/�miƪ�<J��8�e1\9�)b 	+A�>�e��R�^�O���T�?��uS�k>��GȄu��x�m�'E(P���N��V^�3&i�CS��b,�(K���e\1b㼣W��.�4��[\���ׁ��sZq0���=��=p�[��_��xy�_8n�AfKY��8�Q�l�oH۟u�ן���9��*��xf�*+�k��W��jE�#�FgL��$'+.��IH�7����#�p�Hv�H?Ս�\Eˆz����x��Yy �r?������fߕ_��r��F5b��XDZ�N4��w^�5��S������vC�da�9�|Z���;p�J��C��+�l\�O�o����-no��'z䯩'\���yS�i�#���[�Ub�@�'��r!�>f�+���Uj�UK�ۤj�5h\�q���	�ʹe��QG3F��j��"M~ �w�,ӋWg��kx��s>��7�[r�|&h�~��e��v�����L4�S�"����	)ң�v��6��.f�<r�����d����C����X�g�('��lL�pmxGMY�4p{��v8d�,������P�Z�	C��/":(�!憜	H�Uϵ\�Ӵ"
'F|_n���g*�!�<�3�D���Ǌ��.�@�O��_q�8����Z>lz+�xa�e{+0+]�1U?�	�p�ޯD�,�CU߽!V��s�,+������Y	S�}n��!����a�o������<k�`C|����~���{�1*�_�N{{D��� ��HU�-�/�:mt���Pz%�&���y���7��k�?���T~Gsym6^��!	�;T4_ɍ�dg��L�X�dZ�
_�I�[�왮��̈́Q^��(dך:\�����r�hTx��:�L
���|��&(�b�-{v��j �- ����ʎ���<>W[�~c���6 4�P��H��>�DI2mK[ �����c��[=_4��u����M�9iǢ*��q�T�Br��I1iNU��n�K��?�T��[��>;�� u�y��C.\�(���D����t&DO5H�
�;��c��iߍ��7�����g.��t!�ջ'<38��Jw��
heZ���ʾ�rLͧG?�rq6_�c+n:����+���j[?O��r �M,MQ�j�w
c�:�3�WC��o��j-�	#����W���b�����ԬsrI`��:�|��a�%Oh'���3;���`uv�Z�Bm]�Ƕ-����j����R+8��2V��o��/����w����i~�Q�j03�(��;�m�.��7�
Tr��,͉�N�
.CA���pZ��V��O.b~�w΋����/ �z���NwD��� J
����숗f6P���iȡj��+��Ay�F��;y�$搅m���Ы�
�l����,�-�\�961ʏ�=dL�׀Qb{y������HQL�Kj3CwD04�eo:A��+�d�n$�K�5Þ�vni�s7�b`ꌶ��ڼ�¦tw�F�Tb^�d��gy���.1\��a+!pw�q��'��GV�T���ON�۪˟����GS�ex�{�{����f�Wt�0�N��	���SEM{��w(��_��KX%���j�{�<��26oăgp��BK2�G�+�xvZ:��T�BDD�w�X�U�}&m y��Sx�ʩ?�t����.�]�]�&Agr.�&U˸���5Hfm��!�=�+)�a
w��4�/�yo!V�]��L�d�!�@��~Kr���P'�g����}t�	;I{�b�=Ed!��k�.?ӷ�K��0)h�~�j���PW,��p��W�[�^�Bs��6B��R���C�@���û��r��o�X|���K0����"��)o����(M�>��!ږ�\N�o��8۹u�R�m$�����ruZ���m�������;
e'�ڒ���K;��r�o��IGW&��/ �"��O�:S�n9l�\���'�#7U��z3�r:n�%�V�e\�oX���#�L���N�٘�'o"�܆xC7uگ���
32�x�%��Χ�>����Fq|�.�}���w�촿Q.�Ie�(i^مeҬL �<R���b��A�8q8�;?{)1�WӀ�6�� 0K�]��L`�E�3�HR�?������A����>i�gzz[e�N��̈��r�U ��i ���z�������):�<��D��t&t �3�F�(�u�>�L/<���!�7�$�^P�;�@�u����t�#�C̋���Jֹ�z�-�b7Z;��貀���;�#���סw��8i�#�z`�0�q�-|G��ky8�l\}Ã&�2s�ݖs�j��M)����,JE���d���@MRlɝ���������(�@���/x��t��b���4@g�%Z�+v��w�����q�g�Br�+�ͬ�(��2�d�ح�"8tU� H��A/{~�yÚ�l�TK�Up��:Ji܏�����/�y�e�S�(Ϭ*����BN <�T��X�`c��B�%�vyx��(�0ϻ��`�ٺ���0�-4�T�)\�^L�Ͷ�v��nZ�<<4�
Q;ƫ� �
9݊�EJ���*�o3pt�T�LV��htݨ�Ka+&�L��<��ĕ��,m�_�!yb�����pca.�ZJ���;��Č��r^���a���4\2�L��'��Cy8 F��3�_��8U3�w�.j��>�nf���֑Pz�#N�EAm�(��r���M$�S.��%\ޟ98��
!�0ML��r,�f�ﾛT��[�G���U�Y?�"�0x�C2t,=�r�/��We��b�h����B��j��)��k[w�R":�h���Ui�x�㬞����l!�[�r%����#����$�B��P�dKB���I�N2s�q�J�5��_�FA�2l�	�?J��l)_�.4 1�WY�ϑa�v`�)�@�H{8�8�B�����µx�^�	�c<�?K���%D�`��*ڸ��{Q�p|�n0y������j�Uԡ�ݢ_��2��.�+}��8�9K��/�������?�v��{�/eH3���^���=����VA�X�k����ۖ�L�@���M�_��i!I��A7�F���3����eE��w'�T"���X�?,)8����<6��Y�җ�{��t>�.~#����c�tA�(��x��/�ӎ�Sqឃ��u���m��p`�:�[��~�l����X����S��)pI/���AB����8�\$j��6o� �)�X��{B�@yܕ�ս�)��=ú5��A_�"��CX��|�E��J�m|���RlW��~X��t�e����〼&ʿ!������3jjF�=Ieo�&t�푙��V�5iZ$���y-�T�ˠ+�k~{7K�O~d�[���?���j��/� )�����F��dh��'����ץ�|B��)�C�9��2�E���F�M'�<t{��.@zGA.�Ά����M�W��-w<[N5�����Kw�w������% �x��4��@]	�쌂SK�WWk��_���g����u�)�ƍ��\��G�*�h�Z�:����InF��#����B�b`D�#q]#�YN�ud�im��Iֆ����wvۺz�V��ݨ�X�|��(�ோ��h������6~���6#����x� 
|���|���ӭ�$Vٜ�W��B���|�ճ�[ ?!���;�k���|��X�[��3b���lQ�Ҟ e��&�&�&G�A��Y�,`	bw�>%#g~D��^d��3cLk�?��jR�}����@MK�y! �v�1��ȉʎ��U%����50^v.N��y�̦[��(kN4�>hN;��w�ʰI�X0˺���_7.�t;1b�l��ƫ)o$?�Z��p X��!��D@Q$����{,�K�w������i�9�9���Gv[�\����q
�|rX �b>���d�i��]�n&U��+�-݅}f7
�Ҍ��e�4`�F��W��^|��Q�St�x����y�{������q�an~Y��_]��@��v�ӴϾ�Q���
jT"(��3ߛc3D]n���`w�'�Q������QHLdv�M)~l��L�]F���jzDq�a���qܔy��#�B��m����9՘.χ�NA�������f߁�1{��`�S��S�'�;7 k�wI�G��]�P�Op����u�]2�߶�Z�7ȫހ��o7!���P'6�;�Qemx��*�W0�I��A:����0�Z��]x;�;X��?�1S
K�;W/{�B)
;������˷�Q^#��\�c۪i�s�8��Q�QW�V��e�K���r��F�tw�)��R.��"}�1���8�ԗv�z�q���j �4�`�5z��0G�T�ʱ|�b��c��q�X�͖fY�ޙ���Y�sm�ͪ	��eb.�NE�y��(������.`�8*��j��Y������0����UO�O��n���xx�4�A9��1(�~ �8s�2�~�&���h|��q�z�Z��|3a�6�-���d���%�)�k�:����~8{�0%l~��z
��	��X����FDO .s�3+����U���iB��S�a��[փ�7-~�N+M�wb�!K�3��1/$q1Uy��(:�p�by�-�U�]�@Z��L���x�}��)�>ŽO)��#�c�C�_�Ѭ����r��p7z�z%8a!+�Ü�̺=�SżT�9�����ޙ]�Ӥg����4�R��nr=4�C+��IiÁ}IM�)(�k[J驗��$kS�K�%��uR���p�f�M�q��;|+�±��)��@&� �F�~�B�O�>szв��N�/�a��J�����#��/
,����crw�-�cyôr$�e,Mv^��V$�s���g�bj1��F`q�=6+D�R�� z�^N�ٓ�GB�%(�w�d�Q�F񾲠���{�}p-m�ؔ���"���j��3����������
��ha�kS���P�3�%2r�y�2abV���C��}�qߋ�ǎ�}y'Gr�ti�D��r;���9=��f)���$�4�o�?\9Sx�x5�s3�t^���s��j�s{�*
F�hQn-��FLYc����� ����5mrn���Z`v�r�^�&FnN�KCoB-Ј��4�ؓ�������Z5��I����o��P���DΩ4~�����\r�d�w�EqD�:	'�T8L^���n��&�]*�[2���ؕ�Fz�CgE��N�����V��Ҵ#Sq�i�k���Xj�ǣ��̞�!��Q��bzc�<�0����D�G ���T]��h9���SN��+i�ɧ�89�gD��kX�yA���u
U �R�&�.Y]��
���DI��sobE�ic�H�`&��Q'`��O[|�h���|=�y*�w�i;]�aT[<��wC}/B�/���r�F���D��Yc������	�mT�����:j�T�nL�����Z�(�9�K������9�Lxm����֣�����/QJ����B�A�K�@�&�_?B����[�"��t���I�|��Ӆ/�JߎKR��;<+�3��"U�ۨ͆S�*�ԋul�	�oz��-:��q�׿�#�8O�z�Eǯюs��{�c�.�t'Z0�q�+-:���n�����{㿢��v䊗ݡ�1����b�ih�,��67^rɑ�₞�[�W�r��`Zzy>-y�.��9���NZ������?��Ʃ��1]M(�0�Ɵ�������?���b�+�	��g������5'�(��6R�Lc#�L⧁�,P |^���J�-�P!­~D�uO��:&
��H{W��<������<o���_ں�!��'�v�l�x(�ۜ`�
�o~�ǒ��r?�{qg�����[�� �~�h)�{?��0��u6��#9(���'����rz�!�,ڈ3�e�ϰ����U�����3��擘"�*0����9y��y�@�^]��:���ùZ>��O�]�#* H;�jq����BǄf���|6�L�.�`Ձ|ñT�3Y��.���j�v�
�q�9�m�o�E�y6/���,�I��J>�Y|*5��$�.�Aچi�nd�����H�����C��gc4s`0lԲ��v��,h��q��1�_�7�-�I.y�4�0�TQ	n�8S��$`����ưClQw�y��B�/yo�'|�2*�Ma��9�_ᨤ��h�9H� |D�4^e�]���H���Ǖ¬K�y�i���'�D�{�Rw�+�tI	�/�4�r�:�]��X�	5�ҟ�؀pU�s��+H_��֤��y-ƺ:��Sm��wt�(�C7G��pPxaY�Z��3��ʃ�ɿ�x{���|"��;������#����7����o*k��4o3x�0�ʝ�l�"YR£�n� mj��'S�q��/��L��˲Z�\���qNp��!;R��Ⱥ��_
�+��^��1i�#0��v��k�X�'��A����]�n>*"���|���	c'۰�s^��(�Y�r/�K
)�y��f��-�(��1�^�ku�����E�z��������%j�F��6��	��	RPS�E�����w���<I�
Q���Ixr"Ѱ���O+����1U���༥'����7�B� ?(�h����w/L��5�z���!�ם���ƀ��i��������"ۉ!�ڢ����'T�[��*�p�@9.��é8Nm�g��"�>��i�)cG9��Ӱ�:�%ý+�IzĽ�J�+���Nlg��r�����~H?3��q�԰�iM!��3?a��T�L�F�>�t"��[b�2'}�`
�[A("d�n���~��@.�rg{�md�S^���|��B�;����w��(��5