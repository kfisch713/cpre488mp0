XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$i��;`�3W�ׄ�!-"��xh�b�a�c�T�!��Ƚ�����9���>�+��\l�"q��Vs7��$�� dTV�1�kx����L���U7���ir�x�B��C�{���[��K\v�����)��X�R�?�񌣅�$:����(�|Ӆ�.Y!������!�:�B_�I-��T�?n3����>(�qR}�()�ӎ"� ¤i2B��_U��4u�\��8N)Z�3��?j%*�Ӭ���%�<�.�~"�e{>-wY5���!p���Ş�J�k��"�����Z�BTV9|+�O!P�ޙ���ڌ���F�W?,\����Ix���0�L`��X��Y�A���]�Ҥ�V�rt�r�};��ʗ[ W��Hd�!ܪ1�����T䙀�ZG����Q�ʮpd%R����6��y�*z�p�2E
��M
���o��N?���eZ�]�k���#���[���O�YU���SQr�<���D<�/�[f�uۼ�U!`e����O|9��om���u����ڔ2]�ǴPM�� y"23��1��I\;Y�0���7d|&-�����ѧ�2�f�LpO��R������&`�����<��cG_7�bi �1�<�}a���gh��W���[o^f�M����m9k_>�s��n��^:T	�����_�/�>>�i���,��L�tf�X��.�W��}�Yfh�%�`Y�������n��aL�]��RI��d��D�6�f�,�i5����XlxVHYEB    b3c6    25b04�4�);�S-��	�v���|��QYt�t�����I���}Q4��:�L;�vT|��c� ��Z`_]"��*��'���&���里U45RǋG��h�=zx�*�����J�A�h��3p7�m�;!W�g�Ki�L����Y�8�зA�g�u�Lls&R7.Z���ҊP�1�lXv`���`2������<���u�:�������|�}�Z�FHw��`�
?|&ڏD��4��.������0ei�����.@��[��J�¦�GBe���-���� ~tKsyRe��~4������.i)������E�B_�G �' ��p��c
�����:Ե�^$`��,ʝ��~ ���2�EL/���>'Pb�*m6R+#e�1�rP��K��wLI���7�`����v��d�x+��eD�M�x"��7��~�,5�"?xs�����^poގ\��#-h'����e���2���Ӳ:����3c(�I�s'�zSr�tN�`c"�P�����|��´]�ACgP�a�����j#+�V��o��-3g��P�ӭ�V�V%	����0�Qq�aLr����%v�;5�U839�p���V��
7�A��*��������ٳT�rn�\c�i	+���I�Y�쯮��W��}őm���Xc�
��tzd擉��_����a��3�):�_�,D��䨧�9�{�ew�����`Ws�ڨ�dp�ǳ\�������Q��Oa4�hi}�����gV
�X��=�g��BSԾ��8e�p����lX�P����h�eNW�=��F�!A�G�G]g礂̃�,�b�d)2U��#�`�Af����!�j��'国R�۽/��l����MPi�;A_�ۆZU#�ç�D����eB�/k�]l�,�`2���-5V�	ن�(=�
�0���#�2�l�2P>��܇ߥ|���B@	�G׸��ܰ=���e�O�(��-��˽%��q?G�!�ԢLD���'>�n-����,F=�b%�朚U�����]�i3"�<�v�Z`5�������q%m����\��)/4�]���W60��}hg�Wδ[�aWb����[#�Z��7	^�P�+�i����7n@������^(�|�YP�����OV�n3֧�����H���Nf�&��7�Ɂ5�"����9oy+,D���H�S��	�>���L��w� ���1�����7��=�W����
A�x+T'�
��QppH�p;�(��Pw���k���B��ȃ�Z�e�-��ҵF�2!G�"Z��ƚ.1���Bk �A��aH��{<㚮�וjj�)X��cZ��ɲ�p�������L��!�,�2z+<�I��+�(�R[��]:��&�F ]N�8�2m'����p̓�h����A~���TIX��o\s������zLU���(�i8��e��ʠQ���u$�V˜9���ي� ��q�
B�.V`h.Sʏ��;Q�ڤ�y4gYb��3Ѡs4��@�d��3�!2��ڎKW��a�~�KF;��
�����)��΅_)�L�D�&␫��BH+L�A�	L���}�F���؇�%��%��
��J� zw,������!I����9����,���i}\z�T��2h?�Rå����DTKwAu��9)�\�Jo'���e�>�~kJeC^}~��$/# 1I�$���rl�x���j��G䬙Uu���b���������V+��ш���r+\)�1 �Ķ������Τ)[h��v�ZN������CV�f�Q���"7HJ�|#���+��c�?�J��-�UtP�Y��L0#(5Y���ҘL]e�NU��0��$p���)���S�2�|����f5��4بgt-5��9Zl�>7f8�e���v�g�H�	r��o��#�sӟ�Lj��ɰ[pJ4
r�DS�y7�[n�^�n����gL�n������1$9ܬ�7t�rRK���[濁2��YĲH[j(y%����b%��Գ�׏[�i<¾�g/~��R۱��U�]��~r�a�N^�Me�)T��&uj*r�eI�C����2v�f�m�8���Ӛ��f��)[i�1����@ ��uEWs<����ąlqowtNžL�!F�ޓ��m�St�Ú��=E(�Ƴux���ۣ�c=E~�� ���6�\MT���ЃZ�ǎ����9>��A�x/;��t�2�.)l�����|Y�%o�캱�B�'i}���)"_o�g戹�����@�j��Fˋ��g�ڎW�Y�ZLHn�����wk˾�߇~\I�ö���+��ni]�aY;Ń��_�� L�1]k1T~.���:y�
��$�l	��5a>�� JAƩbM2�����W�lJZN�w?�g���k�@}�x����6��Kƨ�_��j��v�
YiE'���q���<C@�7��X=]+aDdȺ��R��eYI��q���J�t��H���-��g���V�������2ҩ	����˥��G3�����-�b+ �b�VmO��"�t��5=y��K
Kt��2-`C�m��'��ٶƺ��Ji��#ʏ�9�&�s	O5�.���%���������BU���y�p֍��jȾX>aq0���C֯"��n��j����,����28�R�HX4ȿ.�t��� ��sdx���C)ٟ��߸o].^ڤ#��sC��$LV��C�Uc��Hjg�C"'K�"�ʤM���{>��JK�QgɄ�qΦ�I��Z�c;Ȁ6kO��^���=H8�~^�*����E��%���_��vp"pe����YUV��h
��1J������0��i; ���7,<�M�ʈ�j����%�#���9	1S]��HX�IZ2TD���
�/�Q�߰s|V(GϞ0J4y����/:�3�uw�<�L!ϕ�V�X#({�U{�`�8�?�������qmh�W����j��Mv��N?���!"�����}���*
���^���C��1�3�	P�Jtݴm��$S��mgX�ՏT�;ӛQΨ8��R�6Q��(��[���=����I`c�}��Jr�؊�ڠL�hڳ�UjſQG����e�f�|�lDe�a��9�V|H��� Gϐ=�.�cc�EzL�m��*я7'l�s+��U2e���Z)�bW_��=H�f�Z�[���pT������W0�����Q�,[���~~?�]���OQW�	Jzֽ$-��\��sA��U]��~�ը'��-;�{���π�~����R��Y�h���@=<�"��(j=��ΩQ���Յ�6f�W��5-�ᙑ��}C3���E�[��|�)�ZM	^�*ϳ�����q$|�#�m_L� ��^S�N"/O�@4)����{E�V�p��0��z���8�����נ0� )]�W"��p+��0��C�c��L�?'�f����:	n�gǠDz>vSZ9�R��/G�;����Ȓjב���`L\�皵�Ը����/�ͣ|�d��A3�5����>I.cp�D$6��}�JDr��ʪ�O٪"^�k�gxɬ3.g��ގ��,9*o�������{��5�ղ��x��I�c�p��1�X!EM��8]t=� e��}ؙ�`"{M�EFLo�(��sq|�.Q�V&V}�oBM��:��@A� 	�lq�Yp�~^��nL�}�d�a�lܠ�C���0:SѪ��SR���Mi����=l2��W	ܑ�ӼJ�_���Lcp�"~��:7'nRmQڒ���(��v�,��WJ'{ѣk7*�� 8�)
�_xO�����4;��1o'?{����!)�2�GFhx��IG;P���3>k�U�$��ԏ%eeٛ�Uϫ�E�l?��?@�w�qRP�
��5d@�B;�-�G����N�e��*z,���"(>#�l�GR�A㷀j�����uMj&BX�Q/��������Aټ�j2C�&��5Te���,����$0sW�0�a��X�D��1~E%Uw�{@�����*�����,��	J�����6V��[�9���o�Q�0�+�Yr�h�P �A:so�S��8(��?]���zH_}�{n�П G�.����h�e �I�����,Vu�w#Lv�>eW��U��1ˊ:4P>�.���|Y't��~s�c2�~!h"J�N�6��Pb
#8t�kl��$B`��Y?�\�=}���Lx@�%�,m3��V�5��e�Cn���=b�5a0�b�.G�֚y�vK����v��ys!;�|�Y��/��x���m�;+�<�)R��6ɳ�?x4�1��\��,8L��{2|�����|@����#���c�_O9�Q=�!jJ�ǘ!űC������f,뉚^^��\�}���Ą��hDη�rm��K��1'.�j��qi��j�d��[�!1J9�{5����^FŮ �k��>����x����� ��T�"~�z~ȳ�4{&�w"֥G��>KwD$ &qʾ Xz,@w]��XJ:�/��w�r��������������v�R���W�y`��H�,2��҉_p[s�ǖ��I%�1Y����[^C~2. �
i����ť��=�D3����b�_���π-��b�����a�\yg�~��	�Ӷ}�X��3u��2������u�V��CS��*9�R���>K�ʤ��PKXy�.ԸFEwv���)/�׏7S�0��%�B�Z�'/��
�+87����YZ#sPEIAޱ��m�X��2{9�oja�3 t����3*��gw�kº�G.��s<z��I��3s���Z��E����Nv]�y���5'}���M>�.��=:` �.��������쟈����(xa��n��T����d�xBR*6�m��( :��Nv�IU43�x�(��ɞ�:r���z��Nϒ���;L"!��Ff_��"��K��V���!te��L�7�W=���=��E�o&�t������O��a�љ�9�30�Ot$���8�m�Yb߰T��a��'9hH�V�Ň�c�i�U,;;��a������E�+�>��Y}g��旛������F�(�����Ob���G̃�V�	�ٗ�!�� ��\e��V��U��K�	��9t��:��Dv��+��iزi��Xő%uUI�^�W7�B�/��/}�Y(S����Ǿ���eaQ�J:5��e�V-�}� {Dy�툂6�����;pQ.�md�hYP1�U�v�|O��%H�'�mC_[��l���x��-�siBe���� ǩ�>�g�VNn�4R���b�  ॓Ő� ���`���身o)e_o�PQ252]`�?��m>�+~qr%����G�&�*��J��� ���ٚ$��J��<����>���@�{�H~~I�� C��M��ۓ+��-�Kǜ@�Ԯ^
-�
��̂2��La���i����zǌW8�i�?^є8[1�w$�e׃��Ei��l�s��Mb�ݬ>7��n`�ʚ�ëך�C	�j*]���{��$�k��GZ�8�N\�9t@��Do�I�tj��4g�SV�j&9�2-�Y���Q]��Ez��ί6�ʼ�^m�m�����B�HMlN#}�3>���52cyU���z��Y5�*��t�I+�Ȧ��S���:sX;���%������\DKw��c���B)��|ht>SͤU*��H�S�bp�-+�[\�bBWU�{6c�)Җ�R�n ��}��S�C/��UK��#	7�f� ��3o���u�hI2�=X���J#'����.��K��Y�)�s �mnd�ڑk������p0ŵ��<��u����b�H!v��� V?S+����_x^��g��|J�\*xQ��sf3=ެ">�g�A��LCDxt	YXf���Zil�����x$�u&�`�E�H���梨-���-�%Vc�"2aUn|]� ���s�|��=�ƽ�Q>H�c��p � H"�ߐ�Õ���<�תZ �2�Δ���niïb�#)�t�ȝ]���&3��q����}J�5�%N�n9�j6��T����1?E|�u�y�AU:E�{ù�%���ѿ�^��d֩���p�I��~�5�B��H�G�m �1�����B��1�nK6�U�8C)���G�t*h��2�w��(�1,a<f�jfe��ρju9 ӊ���>O*(8�.��+}��1�� �dAU�e�� o������`8r������jD�$c����В���n�ͮ��[NRy����X>��wk/��l�L�<>�6�J�I�D ?ܴN��n��M���U���_�}쮡*�0�lcY�%7�"6a�͉�FK�]1(hV�q6rb��՘G�x[Sۯ}�kd�U�}вL��RcOζ|_�m-� ߂��hؐa�ނ| <�gz&�����$(���~��ܣ�G�0AL]Wh�nt���M0�V��˩���H�QqC��!��,���z�����`q~��?M���b*h��s�k�&cҷ�`��P$8�ӽ�i�Nq&t7�� ��%�@5~��d1`�ܴȋ\�C��wG�4��I�[��O�׍*6�?� �~h�ƚӔ�@�Zܫ^����$�K��L:}��E�X'�Ԋޒ� ���O��a��Du�`����l7=���r���a���|+���O��N��(����y�x%6����OhG��u������H��K��:/�ѡp+���:^UW�	��(_D~��e6��<��县�1/�]hҕ������4�I�ӡ��1�d:)I:����{$@k��pqP�{I�.j�*q�L۞��M��k`(և /쮓���O�m�d)�C��9��C�Ul����Ք`��i�K� �[^ՙ��=�-|V?�r��K˱�x����Y���S��a�����S|���lyii�ؼ�6�C���dr���
S�>܎h�]�����
��Vy� �.+i�#)��C�K����d��)�I�q� �p�Ѝ��E��&��E����_1��dg���2��K�w��:��D�Z����!�����'���/�!�$����n�'�O��]��̘�*�{� kv�����K$��@�ۍsR����&O�L��̯6w>��Y�N��Sӥ���<=zA���OJv�jc���DN�t8ԳN_�f�^bk4�V��N�Vr���^ؽ�ߕe�_�6�Uw���o��DG�t�0�p������!E��� �?�Ҁ�-�F�κ��#ç0�Q���	L>+�������8�fv����F����I�6p��D�~ݡ��4b4�>�}�@��u�qH=~��zQEn��q��CF�Zu�]bCTϹ�,UqL
W#2H:B�]��༴��z�h��d�u	�|�u���'\(���<W�[<����Q�5��CX�w� P�e�m{�<���S2�/���E�E���A��2uCo�U�v@�|�x���SQ	��)� ���G�j����_�0���֙V@g���h��8��� .+�Z���b�3Zk}"��H+u�5������}��Jt%���E&���8c%'Q~��H4_�n�;�~�P��P���x
\����]�x� �iK�I��Dg4��5�F�tah)���jv����L$��;�����]�A/e޵$��<;���A,�J`�(���̖E�ӠS�+A��v=Y1�!~'J��vԭm�<h�*{`zd-� �7E�Ò�#\�W."	��YH��_��F�z���9KC�a�`�"z�Q�Oƚ�S���;1{{�~�5����aCb#j3�=�9��I�2�f���	"l`�Fؗ)"0�NA�aԖ���+����N۾g�o�Gr$�S��İ�QA���_�������bb)��I��T��1��>���.����������؆�p)��i��·��4L� �U��Y�zO.R喊����{l����xf����T%܎0B���������Ҟ�~�@�j*�Eˮ5+lb��	��\"����i��o��c�K�<=w�g��k��u#�vO:�Ȧ
�6s(��׈�y[t��}�L�r�g��xHQ{#�U�먍j�����,0�p�
U�&j�7��d�b�+C	8�ZG㓃����wx;�U�Z|�F�"��Co��,�T]���m�-�	�וReF����if\�NZ���A$��A�ܿ��|���JN�AKb�%�n�.��s�*�ZO�-���א�!q����["/�}�]tx�/��*�d������sdxI'�2oO�.���7�\_�(�f5�q
�c�p3ɰ�>����s�_+�	�w�ބ<��u�/_��Rw��}�i�J��0¸���!�k%�b�sZ��)t�U��lQj�{ O����sp���"��p�g	\��I����wQ�z�.�ƅ��`:����j2�<w���� R��*k��_���!+�$>��,UJͱ��Re�Ͼ�����I"�
��s���Q\0z��i"�71K�ݐ���	���F�x-�'F��M������f,�#�j�Ʃ�/줇��ۂw8���.^t�b�k͍mt� ��O�+����h�K�+C{ȁt�g�\:��4ӡ>����"��F�+1��6�XA9?�Uǿ�1`rgQ�q�V�4=0J泋�p�ឞl��kwvuK.N{�Y h�����ʛ����li�!�L�%�$BMUO�.�W\��A��5G�\v���~>/<�#N����H>I����2�l:rl�/���r�,zK�?sp���t�2��9,Z�������Hc"�z2���E���NC�`W0� ���yT%R�&佳��eq$E������"Mxh���G5-]�ԁm�lR��טU��#�&�lZwM}����E�\�=>�2�|4����xZ���FV6�ΐm�,�v�j�G��2�`�2������KxMB#���t������!B�^����h����^�)�1�����1W	�|�^aA��~ϩ��"�`�z,�Νr����q�XH;��O������^Ɨ����K���}?��7@Ԗ�SS�����+(��7��U�$�}��4yW���a���i� �G.5�V��ʢ$D꽰�Knޒ�?}1�65<)5�Ry?����4��;�eOb��U��U9�/z�l�#���%lMl�@���X���~�̑1����Zvb��y\�O䉄�3P�{P�|y//��ZM�X���[��3�_�i���4���]&�4	)�Z!���^�H	l�J�����:˧y@�E�������03��_�Z�YM�Z�o���|ħh���k��[��+$�e��w$�R�Ѩ�0<x�Dä��6	�ُ�i���]��G�e��O��%d�C��6`�)��$��{��_z,����Ɗ������/I��7�h���[^������f����8����kӫL+%�rB̳
	��Pz��M�/�t�"!�Uh�3�>�����/��0�5d���S�Kز;�#�����r ٠���9�Ѯ�)�&BA�