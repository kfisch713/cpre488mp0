XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&}g� �>�+n6vy<��	��0�̼p���2 x��+>U�wQ�SKp�����HUk�
�FU�N
�o$Z#>	�V�bG
�,¼t�޸2�G�drB�<
���e\0̏�� ��(,c6��g)Sh�g�08k���������D��xRY�ۊJ�<��dܨ�2�J�1��룒t~�~�[�>��SU��^ZWa���gV6һ���M�VQR�46�����e�r�I��1KN�(	�Y�ܳ*1�-�`j7���<q����o�J���b��^��7�o�n��Ҳ��#`�
�Dv[�τq_)�y���h��:L�B����t�e�L��˂����fL�>�H���u|�ƐA���$���;M��ރ�N����:�N*�0�n�ǟPll}���+b����G���͆��X1�"�D�ʦ���&X�5�X52��dV�٠vi�5x�,b��z���
(��� �1�� �z1���/�~7�1��e��ϊW0� ��V��sS�C�32P<@x��F����EG�������"� ��2"s3���N�-֦���;MB:~Xtg�Ӂb:Ǯ��I贷��CP��p8��6�|y���E���K�9e��L��Ԩl�g���Y�TAS����ݾ�ߘ��>$B����to�*�\�v�V����?��wI@�m�,آ-�2ɨ �hzO���*kRp��q�F���z�X����^�z?��Q��L,��0��ņ�1�h�:U��[hl�]���XlxVHYEB    95d3    18d0�b�_dc���4�;�xm�	�]��ȍ��@�q��9A���ʬ�|�?\7N|K#�磁 S�����m������j�+q d"aY��?t3c�ZO��6�"{�L'N�Yw���E�;-���R���rs�Hͩ2��3U ��w}�}P�Z5�c).���!f[��H�l�d���>=������0�.��(��%6��G!S��Ƒݏ.�^�hȿ������v��C,cz���܀I_�Z��@�����6�T��i��8�߂��v@J�}�7����Y3R��*ܱ�^���2��z�����7��6q���Q{��y��v�Ѥ0�ѕ0|�/]6��������gg��Be/4�����pB g	#{I�t�20S�i%O�����8E�|nH�����v�EԤ�:?��3tپHu�Y�<�W���_�%��>��Ĉ�l0�1&[���|�&�/��t" *�,\�Bc�u]X�C��ƒ}��3J�����1jY�j
����O3����h�_܂Y�Dx�2���FG��7E����&Q���@����L6���`.	���F�f���fǽu
���h�w� ��Q�Ա�4�'���Ae�C �Ы���{݅T,|��3�1����T���=Sx�/tA�����3��b�֚�#�g\�%��,f,e
�vIm���
_;l��]y[�1f���C/��%z�O��e}�/����:��2�o�Y�):�JE�B%P)�U�dE[88 �業���|�D7;�7�٫�.�9���&w��j+�|)�v��jJ��.���;����f-�ɢp���o��<��滺(��y���!8�$����r��Y�@��eD��.S}{.qHӖ~�`�_���;J����rGg��-a��޵<�1B5�ё�f"_��Q�D����i�nm6)�v}�.����a�j����hI�Xs$�$�{���_��J?�&�	a�~]�����R��26�4X��&ݩU�o��l�
�]�?G#6���F�c��Ia��ճ�3�XM�Q��Z�H%�h �l���ԍ}�$��k3��kn����|��G��U�n}�E�w�|�{ԕK笝惵gr��ѬU��ғ��<��5���BؖX�֛Ԩn�����^�^`1#Dh)*��qDD������iX͡f�Gv�ka��t!���hAe�jf�w WG�m��)�����l�g<�E���ms��AKX@�|?������l���g��I0j(�_����ü*�����d�b"���Cm�u��DB`��&�D����a(��4�>H��.vٹ*v���<�:8SW�ܱ6@��x��P���4�[Qe��b�'����fl��l
�8{�h�����9a{
`��ݪ�>pFR@	�El�)
�WK�5T"�p�?c'��$�7��
F���s���&�����]�o,s4r����g}� %9�A�
y��7�(���旙x}�م���2X @���J�LR���6m����@ Xz���{�*Ӭq#Bk�����1��ϛ�Q�k<�*G�2�}$����/���b�6�
�M�Nb�b+�jт�Ie��w�S�ݦΎ�O�51�d��8l֖��7�S6�)���74��A�ŋ�@XI_u�g�.��/�X�����r%͛E�
�W0���r�1"�I�-��`è1��TW�p&3_��GY�Iry�����iס/H�y<:�K/�	������h���Wb5����3Ǧ���s��p�����Р����W
I=�I�@�$Y�{���j,Ⱥqc6���Ga��9歃��6�,���g��b���wƲ��l �#������4���K��ަ=FAUc�c��ێ�d������9��k���#��]y�+-3xة9W���S�N7$S�l�֣d���D��F��Fǹd�p[ƿ�yI(��0>���4�����Z]��WBZh?����b��C�ܮwZn�m9��KH�(nq�m��ᇸ���`}x�	v^r(x�x�g��s\B��9���}�Uf�]���"Ư����ҡ�iK�ċ�pH�$�7��/6o'���-W��M���^&w����Xr���ᐇ��.�S ��Uַ`���{�I��{>����]��Lb�3����dT軚��G��t��3����hj0���-#��8��������Ob�	����);�~��#S��u��w��C��N{���EA����-��>�ALĕ���`�W�zi+��L��I�Y[�`$�(}���~�ot=戌���2d���"K�A���=��2{ѮB��Y�@�L�N�[���>������³�e-/��uCG�?9#����i�9$V�.���1��aP���CtΦ2��:_H�b�h�6�Ur���%y�� ��(_t���Ƣ����9�A�\\}v
tp�����0�^�V���9�	k��Ƀsϻ�:�7oH�I�	��r��؟�����Y_^r;�ܩ��к��[�<ܕ0�;E#+k�� @
�M&u�{&C�E�B����V�1����e�a�o�1�B_hN�-2��ڮ����5��K���'4��d��G���9��,�q&Рz�Of"�@��T
��kD��i�.s�(
�s��D}��*$��罁�Ӡܐ�p�A�H=�4�N���  �VO8���#e��F��S�y��7xuW ~*,5b�!����&��P|Z��7�3+��o���u)�����`%Wt���"bͷ�h�\'V�:}G��hH����� ��a��c�gj5��'�J[:�읛��7\r�ZJ$�˓��g2év���r'I��I^Q:����
�IW��~�2G\�t"wU�p��AnO�$�Kd1v,�����@W?��q.f�RPh���D0n��+�-.�/Z��1�0 ������Q�m���nh��r4�XZ��(� �o@�բ`���)f��fX��$7���P���1�����H��h՛e��U��12�Hd���;��3*����9mf���X��F5��]U��T7���	�H������T���U�������=�sB����P9����.T��������.O5'������5��]�����w�2�JT<O��Ͼ�����1p�=[��h&}��Xp6�����F�������U��}��U�_�x�夑�J5��UI���M��(�0��aL��*j�W��Ϝ�v��QQ���e��S@Gq�`>�d�,5�f.' �:�u���@�~h�*T���g��;�ѝV��_6��z 6 To�<�-�DI
�NT�`���
�������+U���>j�A�O���|q�N�-�nm�Nu�G��%j%�z��u��PwRU�~l�z���<Bm<�Λ��eM������������x���S�����k[:LB�C콌�}#u͑��h�1����O��d ��mvqw��=y�����~�B��),�wUhx��?s�(ܴP5-��T�Aw��m<���D�P�ʘѯ�=�F���ctȾ΀e��sz��8�,��m9��W�z�i���ҍU���'�3�T"�պ�
S���bSIX��k�~6s��W��,mZ���J��*�<'�&�A��
I����bd,�6�Iz���z7���׵L�2�PâD��J�����@�Ѷ��P5���=�ϗF�#��B��"�9^2Ȯ���0�� x�b/?]������n�e�B��6.���FW��h�Q��[3O�x1�O�[��U���9��v��M�L&T{ѹkϞ�I��f����H��l��#��5
 ˚��M�9��N�gQ4�L��T�N�>{�H���hΝ�S �vAWy��4������'&m8`���p���=M:�|L�ke9�;IGv�{��� v����FѢ�.&gfֹ�A]6�v�b�-$c�)�)�wI4��3ϧ�l?���M(�K�P�\�[)��ye�}�� f��h���D@�����=Eû��n��>��$�_l�g}#u5i�@��Q<��c"��G3{�_!�лݝ88�O���J吺~.{���z_XB���Rp�Ϝ�M�(���������]�^�������N�OX
ü�D�c�v�Eqj��Fz��ca툷���z^un��h��6Z"?����^"�[%�T5����Y�ɸ��u���d�����G0ER�5�1���
�t��)"N�En��J���#$�g��nZ�P ��¹��{�"N�;_�s�]��C% 1p�A��Qh���6)l�+��p|��������9)E`�5\��ﱟn�����l!���H�l����쑂p�cc� �.쐕��ĈQ�v�����q��?&o��"�fgY�`sk~��.��]�]��h�/ڟ"[�/lϚ��ЖDS>h� �o�q!M?{�{�`��}dR�������Ld2dē�8(��f�;�SjX��/(�UBU�Ehʜ���@�gz�n�G��o�؇yL�7rg��Y�'ŭ������W:��"v��r�� ��s������Q�tsm?TY����
1��[^/�.'C�F�5,g*��ɛ����m��S���A,�~�$�I��:l�����㗙����J���F0�X�1�E�yuY��.��e�,NӁ�\gf2;�ޝ������.C�D߼�1Yv�e�$�a�k|>IB�L�ݟc���m�v����r���L�|5�5l-E�qL-�I������u$����䰔'߇A�B�l~�(��T'��f���4�տ�(����s�sS�e*??d�P���摃6����!�UGQ�{������į���'�P�J0�q��ą4Y��,/]Z���f�ׇ
��D���UH!Ew�lf||�q�{���3�t�0L��/��h�~Vw��h��%~K��e�qn1� {�)�0���(�9��������d���#g�A�)��z�]-��	>�S 7U��T�'��ߕ��$�����@�Z�k}&�(����kT0�I�^�[���:ݛS!���Ս5��ɉ��V�yQ<���7�%���ZM�>�{!��Q��lq�j��B�k��D
XH�m�@P����(d尕1#��Yc		�-�����a I݀'T,y�s����P�� 6	�]��h��Mrel�,��s*��<��wpt{P|�	,m��@�D��������04PMTb�Os�#�a͜�H���o�X��P���i?����i��̈���1�|h�1y{G����D�von$�� ���u	�(�T�ӥx1�1�Dy^��g`2V	�C%�Q?x�v�Dh�y��*2b���?�|7P?'8��_�j��K{Q���4r¼�G<]�W�҉<	����3_*ݹ��F�j���3�$�@����Y�y?aC�A#�@@Q��� ɡ�aD��9P/O#����Xֹ�L����["���F��f�9��i%�&�bO8d�1ڍ��&1talbv�i�OН��?3^��$~ϗ8
`�~.���/�`@����H�fnktn����i�nq��"!K�l�&��ߌ�P����:^�G'j������w<�S�Q��ϻ�;?E��&���E>�_ζ|W�q@O�đ*�֜�-�gK�Lt/T�	u	2匒_�g������=/m �b���l?��)m�f�� �S[E�V��K��0z��'�f�bT���w�\$x���ʗ*���#rK%L��jV�����eb{��;�*A���|��v���X�u�|~~��a�dK�� ue��n���"��C��̯5I�GUHC�	��(u�q�p'��{Z��/l����D.tQL˲�����j�r�Ħr�@�0H�y3���e�Q���r�l��L67�5c-�P�4��U���)���iv*�r7"i�x�k�Y�&o�����w�m�ǁ'=�u�I���P��N����Y44�@S5�Z��w<�㘕8�tE�8Mh�ߺ�"�`�����9����;�)��ka�5�襪������0�m:����B��>Z��*~@��R h\�
��J]O��uY�F,"W
1����/���:e����s`�r��˧U��؃1�E�o�v?��/H2���.�eJ�9q%m%T���{��_t���Bi}�W&�%1e�b��uGr��,$0 6[��PR ���"N|Ɍ�Àp��v:���QI"��\�6�n�1��U�����M��7.��u�������+{