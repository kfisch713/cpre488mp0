XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������I��k�娪��qzlRZ{�ܴ%��fo�0���8dz)�("Ӣ�~��V��]$�'��J��FE��/��Q�W��Y �M�Ls����8��M(��æQ�#�2p�׺�\}GpXe{H5�Ϩ���}���ЯF�e�.lW�O>�����Yܿ���Y���Cs��,ׅ��q�%�`�]�z�&��}t35��ט�G��A\��T�%g0f����0&�8z�,�e�K�ȕ'ƷT��5Nu�<4���K&6�V�R�%���!�`�Vg���k�\c�IW�� �4@1��0��aR��Xw��*�/�.��nf|�i{S�[��
���P��<vHn^sk3���!�L�<��7of���~m�	�o���-���XP3�|��0��d��WE���[��	Vm��>m�u��׬��Le�7��jn��6$a�)��0��7�_�֪�V��{ 
KTk���I��j)#�ԃ~j'[��m�˵)��
G.Q�fS�*Ǻ�WB��֊ԥ��k�R��ȍ_�̖��#E3��Gڀmq1���FV�d���1XIKa/����z}bz�J�j�]1rJ����d�o\��beM�a�����"�PTH<
��$L�0n���N-��T薬�Q@��o��=��\��GEe a7��3�Ts�넖2�>'�����K��vS�N�irg#��Gb�����&׺;��������4�BSթ<��Y'���$����
Ub�-
=D%_Lp��.Z$y������RF�9��XlxVHYEB    dd8f    2160o>�)��av��&��)[��C�`-=j��᱙?rZ�}��
�Q��uR��m�4�Fȸ�߲����d��9z!��.@��~�r$_	��X}��VB�N����-Kb�E�)��շ��t,���YJT'E����y��;"��20�c����mA!^V �"�VB��Z�6�3nD�@\�I����ȟ5�1P���G����wdYPw�2l�J_wD`�a<� ���k�1��gޏ5c�v�9.Zs{�IVK�n��KA?R=�@,q�t��=�S�0#oڵD�9(?\u��딳���)�<]OR�@�.G�.L��<y'�"l�<�[�d���
�G:/�#�\��w�M�=��� x�.P��O�l���,<��|:V�j�ɲ����Ǆ�g|9L��[!��S Q%A���J.1���@!n��\j�@�!�h�mH,��Fr��ބ(�^�˝)422�m�l��N+C�E!�u�n��P�Do9�˩n3W~tD�y�C�/{܈�7>�נ�Q�&�FDA��^!/�2	�Q_`�~j���D��#����Cѫ�ÈL���w�zղ���3{9����k.��KG'�ɝ���rm�Q�R�>Rs��h<����Al�Ny��9�E��v�rx�˦VʀLׁ����k�:�i�:���k�b�VN`i������P���:�(�F��e)�����lHL�]�	$xJ�h�L�������D�䖗+X�x#�H	M��2�$�xl8G�O+.�p��y�<Y�"�b�"�xo,�Ʃ�ņ�D߹jX(R�8�0�q�]�P&�� ��P���K��U��9dB~:ɋ{���E�1�Pq���Pܭ�Pc��������X��,0i�vxar�9k���1T��L����6�+�>T`�*�����A�0q�>m�<Q�lV?Qc_1|Y�����@d�w��4%�)oT�wY.�bE#��P0̼�nv��A��~/Y��a�zK��g�o����2��ˍ�����*u$`׎�'�֏
��n�����r `י��"f	1���ٌ�q���8X������ۼn]�����;p���,L�i��v��Y�6q�! �Ÿ9�H ��[׻�.q5�V�3�*w^蠁���������ܢJ�k�rAn#�g*[�0f{��ڣܽ�a�Sf�(�Ka,C���=�ۚ
����L����}M�$��{�]Ʀ7��$�6���'��_v�K%BC����&�5nc����,w��N��t�Z�/U�X�N���凴N�Z����'<.�0�D�ji�ݏ��#�7N�չC>Z�����o#4��zӟεjC�.u��~��%!L���,�
�=��u�T6=��R�M��T��:n�m�A�c�K,� r��M�1+�Q�?�N���� C�X�����7�a�IC<��FMߠ9��Ð�^V{5���rPz�'��P�;��	��v:��csK�-�r]}V���P��9�5��usJ)��kXl�t:v�2�l-K 5��R.=|���(��cFB���@�u�@�O�`�����8�/�#�ȍe�FIDV�}=�o�J���բ�k�tӑZ�0Tn`���P�[}�W��Q�lk��O���Q����ܿ�7�4���d�y�g����H��U��^����n��'C�8#�QҬSi���b�8o:?�������,|5^/�o�CaQ����pth7лE%ڳs��G�=�wQO�qO�m8�{�,β؅�I���T���?d���T���=~h�JB|P�!��dS�iʒ4�@��P+��[���	l�����6?�˿��9�p0!|&xb֑��Z2굹�ƻڭ��޳Q�o[T�����ƌIN�������V�W��qM��P3��p?��r�G�g�l�H��r�[�d���F�������t_��3�s����'شwdr�N����W�'
��!\��_5��<�$3.��t'���&�H4>E��#�S���u�]�[�Cu><w�҄V�ƌ�Tz/�fp��_�[���a}/��<(���hW���z
Y+|1QA���j`_���
�e�I���K���Eim�M4��U1S�7XZC�*R#*� � U��}���e�QC������1�K���G�%��k��|�'!)�3��ς�O+j�����b����k�{xt�_y�$�+8ߊ?����4}�i˸���Č�QxV��W�hak���+��]��۽���1l_��l�s����Y��]؛ 9�V|�_Uj�W���~���	[���!=�Y#�5��ht��#���yW�e�����q9�&$B1��(�{k��N(����y�OU�,��{g
��fqe�X ���q�;�:sJI�>�Lf�.�UO+S���K���
Q;' �"�-��_��>�_��v1��)����Re�u�T��ï������5��q��M<�M1Z��n�U,�����]�g�����P9�
@3^��>����PrK���ZAI�oӬ��a�М���"�eܮ����i'R��l�� ��^�kM�����=%p�v�jy��w�X�g�g2�c=E������W%��ն��CG6:R>��3��A:W��y@k���V8]����g��$z��'zʀ���t	���?��J�S ����Ȟ���7�_ʁ�5�*�[�����ϩr��`�͸Մm\�r�j���u�T���P0ћ.5B�k�*�_lP6J�E�i���:X���n��O��\�����+��t��V*�{��*��3N&�Sd�����t���+T9��\o�h�v�JψJ:�j5���~$k�H�M,���?;�oڨ4ڼ�)̽�N�*�j����c峮&�P�&$��W3�l���+��tL�xr�0��M�6�oZzW�f���f�q���%�:��+,�n�Ң���hlK�X	��H����&|�4�H^F�FCy_3+��e��X���)p0�P���� � V�� �?�	+ip@vn����8U(
 c��٥��^q�!6�-b�-�?�GӬ����ui#��LH
yխ	ɠ�d�z��&�8̝�UL�/Я[���AG�P�`��R��P+��VC�d�A"W*<'�|�w�QX��=[��{��6P�]��@/�4~��r��9��GS�|�%�\�gW��0;�@��t=D�a>��۴��� ��W7O�^s��l�?,�����2���
��,��:9:$�G���<|Ev��M;���"�eC%�(?O9�=�mE����4<��\M~<,�ÿ��]�W!ƺkχ�A�Ap�.9)�����a��eL��m�
!���	�1�
���M����G��Νt�	�10�%)7�zL9!	�ߢ���fݜ�Z��g�q��ۏӁ��FBڶ[|B<��sbӈ2F��-�Ҋ�l5�&�i�J�QD�!nD���L�e������M�s��E���3��XU�G?�MW؛�!�(U��M�S�M�3�줆Ɩ���*�s�u�H�-]�P
�0R$d>	045���aإ�n敼�ZT"� �m��Yс����$i�ddbhX�Z�\���!c4�,I�la.L$��;��z��a�S6WD��|��&�
0�03���fCֆ6˩�a8��§v�9���&7���"��˨�����Di����Wpʡ3)0 �\�}	8J2�-���^�Ԝ�&^��Y�e��?N_MW����_ZU���i�RI�$+[�v:\p�jkRMR���H�����ti4���SC-�s��ѐ��V����-�+��O���{���-w���>��r�sy�FJ�1⎯��`Z�T�6hrw���f��W;s�)����n'�_���/A���o�%a�?!�Sr�����t�V��(SO�����q�����Do�5$(�B�h'����ȵ�iS���.5۶��^S�$*<�È^�ͫ�?�+]����t2A(xDx@�=���aQ7ǚ�����½�I2!��6
~���3�y�$Z��]���JT�.Ӫ���� \��} B��'�0�`�4�<�Φ���'�j�D�[�����&L�&mTP�w�r�ځ=�b��Vzۘq<i�&8���$�I3*�ؖ(p����fֲ�Xۥ\J�y�Y<����Bo720)M�(Pr�DZ�H��{�7X�JNf����0�?��l",����D���5�����-t���*��39W��qߖ(`
?4�;�����l�E���|�p����@l!�G��}��Lu�	/B}Q����P�dU� �R�j���?Jz�I�wEk��m$�	��v듄}΄ �mx*����i�${�_�Q����0!�{o�8��-	i��qg^�eT����šS�n33</��x��|ӥO��ܳ&���4���BN�͵����ʠ�hn@�������_FQŮ�V�"!v�x�})W�����ye��Q @ɬ�N.��#�� }�/.��xI�lzj(6�����/�W��m��>�0&Q%ɯ՛ l��N$n�#�A�,y`����&Ԝ
z,���c�iv��pZ�B��ɟ���-%�hݘ H8��ШZ��3�ٓu&LW��1= ��=P�t�&>K�}�\B3v������9ЎYD-e�LE�<���4޴�r�p�!�����T��	�O<6n�k�f��x�fٹ�z!JP��sl(YRkO��KWİ��ӹ,G�����o��F_���Т��H��0@m��2�c� �6��	;�ǦFF�ug�1[��BW����4�H�g��lw���ӁK�K-'KsO�m`9 �3e���:�qnJ3>9a!��x�2H�2e C����J���k�Ǖ��t��KC(w�6�lE��	�.���������d���o��H'"�4Ǥ�� ��I-�{��� �{H��^�9�[��;��;܆�9H�s�#^�h�p)<�jK��I�ZS�3��\�JF�y\Hnp��݁,�j"��������C?���ҡ�}9��XJ:6�oqqӈvF���I�-�7A�&Tb��W!&�P��v�~�	6룣�+:B\���'��Q����%�	�m#�o�}93Ϥ*�҂���r�6����:@M�u*ZS��+������I
�Gq�E��rF����JN}Pg�cb�qԄ�ﰚ�����IW�-�8�&����$�'�������P��aU����}`k����
j�As���Vb1�8�V� �k^^�4��pR�}�D�2�	���Lp�
�|�JU�G�-���G$��L��5���qCը�C=4�9Xڮ�pV4%�xF��*�՜�H���'#d���#�wE>@���1��J�\�zG��ī�g0Fڋ�)uͪ����Ւ��꾯�e�sCd^�x4�ӵE��*P�	��G~.��e�6�!V]v��<X�����4�0�q����彫A�|�]����"�t��Y^ڭ� �������b�Y�����\`뛷�=ݢ�|��D�Q(���0Ӗ@�y�{4�]�NXo����cż�G7�B��|Yi8y^OQP�v� �.k�y�A���N���|�{��X�۸����*��4�
���Po���,���Μ�MZ��Z��t�w2%Cg��Y���
�,+���g ����0!��՞ <h�����!�h�j��}�n���G�SI����W)���Y��+.T�it�JI����`�mzã,4�� �2��(�ە��g�Q銜�l�T�X]�+H���8m��O��\��pM��\�x�M�=p~��^5��ܐ�z%��U��
��?	H0�9���<��Y��=��q���[5`XO+�ܣ7����c�~�Mܮ`�u�`�Vc|�j�'164�<uZq��U�������?�(�F���:�7l6�6�[�hdO�7[s�����ajwɸW]fSa����U�L�c�-�{�p�R��"��V����H�E&f�j����EԾO�d��D%�PJ�eS:U�����e4�"d�����GH��>�-����JnXkQgjn�S�M=�VsҠ�������E�2>h��3�r�����g�����dq������d}k��(G1@��"��1E�8�� ��6�W<n��]j��4n賿�����4{{wύ�T�Lol�;%�������H�v�e�ѭ	� ~�p�P^Җ't�0��x%�Vj�)��\%��ȧ���ɮ�^�4�<�s/x0םuM ,��^�<e��"$[طK6D�Sg�� N<�M���g���"ˬ��w���,�sj8�p���8���n�pz�Pcݭ(4$[�}�+�����L��	���I �a,�����0I���7����$İ��}���B6}u���A�B��h�ҟY�d9���9�#[�.��/b>;�8a^��i���
/$ݜM��x{���3�|J��0��I�s0��-��X{�s�e�@���7��27��m�$i`����^l�|�#d(�B���9�e��3�}�O�T	~�l���O����S�J/֓+M��[5Y� �ʐ_����a�Yj0v��x�E���_Wi�XoC�$ҳ�5��#�d�NՓ����[�ǳ� B�������H�G�LڕǷ3Qv�R�%�9-�o�Glb38�s�Y�	rАNh���}�
���k�/u�	�jlr��s�M�� ����Ǟ�Y��r���>3V�c" �'�R��~R����k�fb[RtK:��9!B�����Rv��;:DcްdW��
`�ćD��pL�E`A��0X�F�YIE��-n�f���LK�VB�f~Q�[��(�NnͿ�"��d�k�D-�rE.�殺ʹ�b<�R�@��*-�ATی�6f���׎��Iřp��]�#�l�@�[Vԭ8FI�R �E��D�JI͊JhT��
"��=��!&r�pC���e�>زG�O�NY^���!ތ0E�K�%�i���/�����V5Ѳ	y�7����5�%��n,��?��n���n+#�VUJ7MOhً�O��Б̓��Y��+�-;�-'K*�0�|�O<�o	�┞:����l�-;�f
U�KyD�_�v}/�o����̊�tʤ������%�b|6-��
M�鴋O_�����y/�F���!g yƙ{$������Qmt��6��K�q�z�]�[ٛ������F��W�<LK�e�u��Fٱ��5���x�D�~4�W '-k�A��=���{;z%�,��DM�5�蜀wv�%C���e:�٭��fd;Â����k}M��uW�x0��M\7��&]*�z^xR<����*��M�3�W�G�2����8��׺���0�d!	��C�[;+�� G,5�dy��̿;�3�
#���{����:���-h��)k��.�-�������S*���C5b�J�ͫo�s!�+0���=��]N0�c.h;����BG'�_}/�g�&[ȣ��m^���3BOĆ[����g�M	���(��S:�%���3� ��m�Ƽ�lC}����-��i�[�`�MQ�6(4kw��R^��{�=3#)��`t4ف�/V�޿��7�* i��8�+b�r�H������m�φ�20�Y�I3p���,�iDʡ�N�- �쭙��y`$ݘ��a�S����˖=�����F����j��P���;�ia��Q���-���ٸ��X�XCz�"��*
���>;�j\u�K������%z1�d~�PD��7�ܙ��Ir�%����d��� $ 1�����l�U��::h��(b
�F����}|��NO�O/#���8{K5��nw?\;?W�]��"m[��W�h�]��y��Ѳ��4�H��_fU�rW&ͪrtk2t� ֓��ͱ�9�!~�}��bs�.��Nn�x��S,��X�L{�eE&Sٳqǚ>�`1A�ǵ &��Y�r�;�<H�'x�p
�`C�QfΪƟ��������K҈�xY��CS��33x�z�����^������:�Tё�qM	P���V༙�f�ζ@��t��)x;���N#�HKX��ʯ��"@�)Gq[�E��@��VKLB����k{0�B]ÃA�H��1�U4��Ę5T�5�@
8�ݮh�7���DL.b���1��v�`m�q+�מC�v���*K2���@��O����2I�����B
^mW�&,zH.���N.*9�#�ĪD��b��F�Dp����65A�ɗ��l4_t����|0�(ߢ~����	Pʝ����B?\�t��/:W���n@�~|~�h	�ht�8�d@3�g��s"|Q)=��h4 ��J�����;X�a|<�-�~U�s u��r��I��m�[�B�R�(1�D֜�\a�`i��M����T&����m�oQqHF��d	�?$ɯ��-�0�[:29��i��_K�	�lP���pv�>��Zd]����;�