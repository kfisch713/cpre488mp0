XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���-Ҏ�'W���j���_����o�s���.*�N�������-��OY<J�Vn(&�f_�q<�L߻�-d�)wc��6�M�C����=~涔ӧS�=��|��PC��5�y^z%ĺ������;���F0iG�-um��ŵ�����[���eD��ODmUW�0�4SfF̼�y{:,��ڂ�Z��|�d���K��
���l���T9#r!�sh�du���%EN���!�;��\�{X3�E�,�����t}�><�2�vd����E�֜̿0}�?
I���X-RBXA`��E�w�
O�L�;O���p��@�R�??9+�v��q��u�9AᎣ��y����_
K_���m����O'�q�Y�oD�)�Vn�U�p����	<�j+�PH;�S�����"���W͊�*Λ��z*(�?�c;�ǘ�?��XK6��b���"����0�#-�u�����Q󖥻�F���[%��c��T���6�H�󺉒�H��\�ޗ=�i;��Uc��f66�3����.P0~:C9�b�5�<^_<��G��)e�?G�Ak%���,+���(h[,��i`�!�{�y��)M"G��w�w%�b=�=n*C?�[�tIٴ���l�/� ��O7\m}e��]�	7X��}� ���,,J/lUi�U*�=��IO
*@$�1T�Sh��c�;=.Q.C�ə]ٿ��M	��v>_��;Nbgq��7^o}�Fa�˦����dXlxVHYEB    6346    17903��RV��w<�&)�d&$��ݚK��D�
�x�(j;-nX�Z��xJϩ[=��v�V$d���pL�s�UOY�L�$\�`lA' L]sy,o�[Ɖvu��O*�y*�ᚋ|����9�Ri�6o_0�<n>��8�f/�'�y�˶y49Q������'E[6}p�=]82���c���H k�gK����/Φk��+=q"�C�*#Z͇E�w�<QbQ_��ȕLU�>��e�Pb꧄��I�q`i��-#S�#�X����BƢ��,)���/���-���v��g|p ��A�AZ����J�H	߷/x#N���ZnU��c��# �r M���.* ��f&��7������ U�y���Pņtؾ�Ĕ�k 9s��A����\+K��F����n�n9�S<�w�(}���r�ƃ��E��h���d��y?뀅� R*�Ȕݐ�+o�x!2�ޮiS�ٗ����.��+LYC���ws��j��!d��3���M��I�� ����Ϻ�W��J-�h/�l�6���_T��A�53�"��;�90����щ��I�{j�%C���&���t�t��-�.RG�eφ����-���=��� ]�@����J���j�閈�8lr[ �x����)_�3�'���W�
%BY�TT�w���X`���3�6[?����Y�~��WR���1�K|d.��[;����|��E1���e����DymQ)����zn���qL�N�TM�9�K&ڭ��o��"�R ����x��=��0�ΤW���<R����Z�@��Ǡ9����+w���>~^��{Iڗ�\4������>��rdf5�è3J��/?T*)H�y�u�����wǉ�^���n�>l��
��E ����~*Ԍ��x����-�W�螇��f+�ܔv�v��RA��'�Y��ܟ=��y�~��Q[����m�)�;O�k�8l��ݶ����ь*�hS�����g�i󈫥S>�
��(�YB�L�����n�Lx�SlûY>�r�dK��N�c�%tv�!��RS/�"C0�G��ְ{f��J�)��\�և'� �0"L��S�Ѻm�n����(Y��p��9ò�g!��츺��Fw[1�b9N�X��'��i�&Q`|�~/�i�C<��,#2!+4<%�	�-�$,�4c�R(S�c1j�|�g���A��Y�F��ƶ%�7L�ZN-�����uZ�����1��QD�ӟ�h�y�਀lȨ2����A%J L��#�L��e^��};+���4?�? _ˉ���/L'�K�r�U����Z�Ox0����Vi`AY�@$/+oNVį�n�ϸ�`��0i~Q3�Э��o�F�׾.Y���J���nM����#�����\�؍��~�����O�l���'��]�d���Ak������$7S����3��d�h�hi��!n��6c�x*ɛ'��n������������>D�6��՝�:;�l��^�=� ��gL�'�}���-KPВˋ��.z�+ pr�<`Z�a��
�Ʒ
�ó<�E ��51s�1�N�Ztx�=�̆�1G�9���W���`��؞u��HNf�X�4���q�1�`�٦4������5,;d.��)��omH!�Ua���E����vy[���I��}rE�/�$i������L�׊�������4��"��Y�y�,�W��#K�qB�\߲�E?�B��?!�"~�3�8[$�ﲓ��	ފ�e�l�"AoCjj�d̥����I ��*P��$R�Y10�����iF1M����u��\�K�(�~J����͚�~�$!~��u�a ]�`���і���xF����w1�&^Z�r�s����6|�.�i�Z�Hfo�qq�G��BRP�;dzXǴ(��*gBRw�)A��!䛤A��hG�u�n�t�pt��Hi�X�����w�5�͝�� �&\�BF�1Z�����,�na�O2y�r�"��Ar�����Q��&� ԥ�p­�&gj�;�4�j,��K�=���،l��k~ԷH�gk�TUx���ʐ�9�|���s��q��w챇��#�"�G3�6J:�0яע���El�K�D��X�X5o[�ӝ����d�DN�1���!h�o�D� a�8dp��(E���:z��� ��E�s`���*�D3^ij�%Τ�3�P�]��˙���BA�U�a����?a�):?fsTZ����.��Uy���n+J:)4��I�� ѯ�&�_*��*P�U��W	� #偯VpVJh�'k\o��W� �r�4&�ɛ��@P�u?'�t*��pE��[��=W.�O�����^Sod=�]�?�T�����#¦��4��>�{Տ	��5����\< ͫ�i�@�s��3�1�/�ګ�h��`݀�6u����Z�Q0����#�m1�[o���y�z�:���q9+��K�7݅K�'
o���d���������^$tݦ�/+9�[a�
1��fJm���n���!�Fg�����KnrL^�p��!fKC5�>�|6Ww�U�'��|���
�8���P$ۋ�6�W"���ɃX~d��"���q�cC��Z��5j4���|0�#`��1i�S������p��DR�G8hE��>9:f�L�
$kߚ�E����t��
�F�d�]�X��d-����]iYe<�;7��O�}�6*�m��t3�,8y�_��!)T�6D���I9Z�?���g9[5^���h�!�P�"���n�B	ͼ�j��_N����!g��'�f�|H��BX��a��	)�"�|QNVJ���ch7��ߋ�6���vn[����;x:M	R���Ƣ�5P���l+`�X�ɮ�Ex�^d���a.��P�U�c�VS�_���u�JŤڶn���Jp�ļ�1�3G�����G�&�f���Tג�"X����昅�x�2ĥ*⤊��'��eB?
O��b:�_��
@[���;����&7����G��I�V��_��%��h@�2n�JW����S)s!H��� �S�D	$,�|�ޯC툰��~�1]q������ǹp�5u��A�! ��M_wu�����%m"��)\���=�'��'�r|��h�!���ez0OZ4�$x�c>���֠�0Q�z`}��Ny����U�H&
L� �K�#	v�Oo%�����I1>L�l�ӰGc�7W�F|�.�
O�aE�a��̾91�e�����,��iy}�e��]���CK�L��e���E�g�IK�T�aH\�޽��grX	�r�~���Z��M'�Tc�}�|�^@��v/��̩���_L� ���a�'�|��X\ X�5bJ=�R���2B���Tq��ZJL�!?ӯļ�Jv�8>��ͪ7vEH�2���
�X%��S��v� �i��tL��ObU�墍i,��U;��̇Ȟ��#4ǈ~$rd����cG���5�c{v�47�Y�A*y�wK�uR�:��%�->A�]6���q�Q�m*ՙ�D���dL'��:�l.�E�� �G�C.�-AMΤ;�mP�2H�	hD�q���olKv����q?�զ��`#�DӋI�u@�*ASb�ǯ΀Wr��73�|�ja������Q�2D争g�;L����I�p�#t�T3h�u)���2�+J/#����X�{�h#���]Z�ǚY9����~V�Ā#�O݌��U�<w�9��|�e��?oA��9�އr�K:0��`�å�~���[d�ɷ�v	�wr�蕋���S�:�%�$���An�thމŇ�$
)nXD�V�K�[Z��2����~6s�.��v�Z<�3|�C��[:D��X�E���F���ũ3w	S¤*�����
�lZLK?�<*��Lм��5�����*��A��ޟ݂����| ,Hü6�y� "d�<DS��ū��xcD��>i��{�I�,=)����]��T56����.q�<�5�x_���s��
��0���O�}�,ua�Z>����fNN�k�t�}4���t����eZ���N y�xw.2�C����l�`j�P���6���#\�D���7�H��/�!{����K�K���̀�Vǫ?��,�,|�Ng�T�:s������y��s�e�`�*E$�!M��
�mT;\���D��S�5�Ih���KS�a	s�����ISG�o���C�S2tا�\����&]t����A&�q�]`�c%09~� �^��;�PD/����]�ߤl ��\�*�+��N�^ �-j���BX�*F��Z����O�/jV�[���볤�@p�יN��d���/���6�3�)�Z[j�� g���o������sܫ3ү�C�k=����b�����d^��-?(����ޛ��p$m��ެwΎ��U��Ё��IG�g���F�R��d�U���7���'	�X�8HrLi2�A���KG h��w?�֕�m�����^�6���V�%
H��n?��UO�q��J���/���Qvi�a��¼s�V'k	�6��8!i�)�O\d�׵9&�L ÏU�rM-s�#];ǆ^gWE�W��٩����AQ,*)�6>�����+z��~'���fj(�&T�c �,�����`*vӊ���]�4V����nQ/�3��6�[Z9�({툸�>-`W�W�tT"_�}n(�k���Yo*�n�	�,{����AF�ZD烮7�Jl�����EN0���q�ۗ׏�0�ëj�x��T���d聡������)`+����֕�v�^=�Jo���&���ͣ�����rPW�#�иe��$|���ш5�աW-�}D�ׂ9&*�}"�6d��Bg�[���@�B���M�kI._vۗxF�\�\ggS���-P/z6#KzOc
BH��s�rXx�(�h��͹:~��0cU�������L������ۥ�4�U�6!�3Dq�<�̓fԨ8y��N�������U��ج"z�	B�6��eǍ^9k�3PH� �n'�p�|�(�%�u)}��ZU�y����y�C�Ս�{R���?���Z&�Ȥ�{m�㍢N�N��dp��O�;De���{�¿�
`7UR�y9�����-'/�w�vq��W̯���	H�wF���9�**�u����K��7��z���zM�~v>��9����4��p��_����BZc��)U���~~�j-N��D�*�t�]&\v�Uۀw�AR�u���˰���R�B�[b~�d�V:�x������OP����v�u2�{J����/I$$�W��W)0�g���Dҽ�k|��u�� �7�VaKqeK�.x�o�X)�'��+���u_��Y�m���yq����	K>����5�_d�E�ݍ7N�Ы9��	}���|g�b-�]݀ἀ�L�����g�e�#bR�1�?9���ő�a�ˇc�F�si�O�,�_U�<���wj���G�Gp+g�O[�)�8q�q	����a�O�!3�����ja���g~����ڥelS���Yw�q��Z�B�
J$~"2H^�y�[����~8����W�ؔ��P�lo4	�����I*��F��O�)�v����wL�]��j,�?	�` �@��UZeZ!�(v�������������e�+��S9�J}TH��:�קtM��nN�N�~å!����]�:lU������Wu���$5��ʒ-�'�[��µ�T��l�����y�<�������hS���[Z�<�g��z(2�2nCkN��Zv�ߜ���V�q��X�:��j�K�51�����mļL�W��qkm��ۃ\�Y�����
�?eZ"Q�&S� F�$�=MJ�;�B��٩��;t2dآժ������"��