XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����WR���Մ�����K�'�i�¢�mX����������}2�:Z�U�{�=�E�ߌ���:[��j��?�@��;�}�2kڍ�ݎ���Q`��� 縟��ܫ���)�:s��Jp���PX���&���R�G �"k ���BB��.L�k��U�x�ɗS�'�8�e���1mF�_��y.s_�-.�c���w��	G~�g��ұz����G�L�괗���⫻������At��}�i�C�Y����͝j\g'��Q����P�i;�D��͕*�"`�GX�$�t�ZR������ӨIŏ&�3��N�-[��:�V@%�:;��q��,ㆣ �fl�Kp�Z�YZv����fɆL{���,��O����������@�4�i���g�G��> {�3	4G����&%�K�������\�,!m�Vh�(=���e�?���n�>���Ty�ޒ8�z>�Y�c�DNl`�� �r
drn�h�:�9��0 cQ[�I׏S^l�ܑ�z�	DM=}�qº�X��"øFኆ	���k��Tp��$`*J�.D�ټi��� |�)W���%��[�l����
T��l-9y���wr��5��vh�x!�t�R���p��SEeH�\W��?�n�,�:�&o�����/�e�����U�$�=xL���m���QtX�fF�ϛV�~}�,���r��i�	��&g����ǔ\[T���;�l:Μ��t=��Vr��gwB�AJXlxVHYEB    95d3    18d0Ƽ�l��\�ah�a�����/
:{&�z�rG��s��ލQ_bb��--o{���ɏ��_P��r�2�u9��{��ɉ�b(6�ʭ�d�k���Y	�	�������ںPSZ)[=�	kV1_%>i2�N�%vH഼5/�������9z�0I�C�́��;S:�A�^Z�5���i����o`a����n����ed���K��+�51Rv#kbwtD��E�.���
�i=��2�gO�Km,�HϗaL���N�ߋ��AO ��������L�g���X����)z�)�
�<���,�)���Xyq�r�����
'䠉icL+���[wX�բ ���uI�i�Q��4x��p�탙� P�>���~�#p����4r3l��ER V�,v����W���m@5�#�Ůu�������*e��]��Zޚ���Z E\�7,�^�ק�A{9�?�'e�II�&$�=���`��Ǉ���ӑmn�@&��n��R+�3�i�B��"������u��޹����ofC+��R'.iм��M	���}n�n6T�;u0��q {f��L� E�M��ȧ.(���CkD�|}[b ᖎ�j���v����|Y�Q�����)����nᆀ[������!l�� Lsˋc���P�.��,���[���̣ا�7B�ݘ���F`�)�1�H�(�3xK�)��5����C17�忦7����䀗�~{��h���Ly'8��z�{2�(�W����ix2+�5H������rY%6��P�~�ŞhKh�!��F{��DS�a��}.���o5uR�|\��7�&����Q�G\��5�	X�{к�q�����;����ei��z,.�yUq�&r�]Dc|�0�sR�ƍ���7���(���xf�H��-Lh��s�l�]�:�u����z��
 {��)���O�&A���@Iڠ&\o[Vԍ�#��Z0�4�~l�%t��君�h<c����*�Q�p��4n5Ru���
:����`�D��7���#��Z��}�-0qľ���i_�<:�DP'��H�1����J����}I��"}�U��H{�'�-K��*]�EZB�il����O(h-�Yq�yZ��E^W�+��`)�?�3P���H�Yx�o/bKc��Y�OP��P��3�{�b��a�^�/ �m�h�yeo՚<+�O3����}G�`(9.�|����X����n����` ��G� �x�L~��-�V̚'�K���{�`0�S�� k��"�3�	�N���}�2����3ŨՈ�1��X��]wo7��C�<[Z&�~��n����FW�X; A���k�d�/�i����Ҳ�y�������qج����ʣ$-	�9W��[&�e�z���*g58L{����!K���Ap7�3���F����z�L�x^,�$Ki2=���<��Ԥ!Y�8���q��lxB[ �`Cy�ǆ���"pܢ�G��*d���<N�:����4�ȃ?���J��Q��V�r�F]#��~��e2{ߎd�>PE
��9.].����Y|��i>����L)���ڤ�_��+f?�.+Ҥ��.1;��1lwE3�:ȓ��D 1�1[��M��q�pW�rM-_P01�B��i2 ��~2�@6����  {˚AZ�?H�R^�����yЏy}�Ӯ�����A�!�w���6��<�}��(Wђ;�YtϪh���<���hv��켪�ĭ��
/ߡ�2�\���@�| ���sG���dM���ķ��*�����
Ee�SA#�o�Fi��TA9��_E�*&���IW{�Eo�6[>L�ˢ�f����1���h����$Ɩ���C�S�&���:͋�jGq?���Z��,��*Y`<��P~����JrϲVd���jp1jk��9��.;��{�O�5|@C[����'Zg/��q0�c�I9Y�Ss�yS�4^!-Y�W�05�Z�i��g��Z�^᫟a
�
�!�����CRG���B�E�ʵy�$liXyƼ�Ʌ\�se@��)�9����K���mf`��
9��ؑ]-4�a�M�1F����� �� � ��)
��ӓ�R
�X,5����g��+����WXId�LԪ�9��Ppu��<����-�>&y��Z�$ Tk9m���ܥ\�%�K�����〣��ͫ/�R<%���m�gh:�!�UR3I!@���'u�Qkj��a*��B���{�WyQ�|����(И��<���}�9%k�3���m�D���!�=%����1��;lo����龏k妝�����j�v0�63���ta�A��-��M�0���⫁���*��l�N���˥�2�9�~����d�x0:�<"c���OgK����r,
{M�IC��$�a��_b�����_4����8:U��#'Ef �gś�v}"����O�ͱ�;Kˣ��rX����F�O��*8#���D���B�oÂ�j�[�SE� lѢ��d9�<P������㭄	eh����Ή4��0^S�TښN�av %>�GM�L%�ZB��:5[ND:��t�'+Dr���*��7�գiYѸ��G9��. ��)�l�[���[�}::�p����@Bi��4�����WZ�k���l�L�ef ڃ�m}Ր�AN8����̂�-�Z6{@G^�uWC���8fuV�d��/��ߞ������&f�o{�w˛E	EJ��]�/e�ң_����l�o�ۭs�(�Ĭ�wUA� kC*��{\������U�^|��Y����;�K����X9��*�g��f���W��e�c䵄s~����bȺ�ǑH��9� �J`��%�R��.C\PT��~�A�:&b���`L����Ibh�K˼*8��s=��E =S�E¢���Bߣ'�v&����Qwפv�H5��EJ��`s/���U�J*v�T�D���U~!��)X��2vFS���g�('ŐI͇�Wg��s�Xf����ƾ�{5϶���Ηn&C1���]��>
�P��s������-��<��c�m!�V+��e�ֿ�p�K����<@�YM�+|�ٖ�ڡq�l��<܆M.|��:����^�y
�7P{Vs��T�ژ��w���~���Kc;�$&��`�2�޽��N���mۓV�
�b��A����Ow#��i6 �@��i{/�xG��"}�K뉫@� �^�G�
�H��G��W��%�I��8W�G� ���Y<u��WOZ�;�V���C�na�P�p�j9�3gj���Uh33�����-b
p�z�$�0x��iiL׶�������&̪�j��&`۲�%��v������{�>�Y.n|��MS��� /"~1�n`7���j+q�2&A�]�f�� ;�[G�'Y��kb\��>�Z$�e�a��H��D%������l<+.6�,U�U:�͛�A������p��&UwU0c���z��`M~�L���{/�/:��Ёe�K�FS�Y'�/�F�b��w��X�5Z<S�z����q����2O<���+�i7�E��oD	늡�J�q�7��3����Q�������M���&K���=�?��4"��a=f����
ŉ��Gl�7�g���=<?�Au�|[�Z��������P7Y�f^P��q41�	�
ǐlVk�t����툩�M8�	I#)��\�Y�N�t��r�cZ�x^��@�yz�	���5�ȏ��&ٻ��%y��wU���jߔ_7����ҩ����}�ߏ�@ �����8R3㙳������~tr`�}�?�C�0pf�Y}G\�»Y�W��]x��R'�뉃�^u�j1��#د�Ǝ�OU>�&����l�\��[����������
ɀ�i�b���������f4��p�뵡>hWEc�a�i�����`�s��۱P��9;K�&c�hnRE76��ӡ��Xz����RkJSg�#P#�>�|��b:�UϢW��6�ɣ����
%�E{9��jݎ��*���2LZ����d5ˠ��)X�#[���� eFu?9�ɗv���y�l��!�`|l����9�5�=#~>�:	�X����\ýc�|+���mK�u}(��g��1�zI�]P������c�ҥ�,cF.qܚ� �v�������/F?��.4��\�:Z`���u�{�Zw�x˒�z�A�;�H�P�͒Y08�움Rh�d�\bU3�+�V}�y�͜Wj|�'��d�I�ܼ��0#'$���Cy�ob2�gVث@S�O���s��]�Bd�2�y����U�Ӊp�a΀ط��m�p�1��|��6u�#VM�����e����E�_҈t<�)C>�����{Nn�L@|��1�PT�?6|�6h4���M6ǚ��,�Y�Y���%����a��L6��m�ʹ��R@K��z�8`X��JkE�� d�ɘ1��\��S'�I����Q@-Vf�0d��o��x��S��-����3>Ĭ�'+�'<�3��'��R#��G�����&+t�wȠ}�iᗢ�M�_D����+j��ɟW�>$X��;��6�(I�u���:�*�_����Yi�Ύ�v����Y/A�XY�z���X��=ɰ�J��0��Ś{R�$�+�כ�r?����.W!tҁ�"=:0�\G���+�q�	 �oIݕ�4���s7���yϤ-A�c/�<�Ϊ�u��W�v���2�B�Eֽ�D�^#��8��g�z�x�"g����M�NkD
�t��?�JT�'��QC�� �cDH�	�zh�|��>�X��V�|��_��,��(3���E��<�E�u����F�E8�P2����� ���y�!�e��s۲g�ۢ�C@�Wi�Zy�J/�4��BӄtZ����Z��=Y�A��l��t��cQKg�&��e1E�΍M
�ȫ�}��<N��΀��᪟���d͍���Ap�!C�͢"�-k�Z�3�Q\(�}��>�|��^[���0�3?ֱ��PR�K� ��_�Z�L�d�� t��v�@���(K�����ߑj�\Ը��93�>�(��@ok����9U�T�!�
#QQ�|�ܾ��EY2G��~+�DAιW����	D��̴�"�ԡ�5:��'�.�D���d�iX�X�d9JD��+�WIi̿�9�����Ԋ���3����j���ʚC#E,��su3��z�����}��?�Ǡg�
�v�b�?04��ø�
�'AC�P3�)p  �"� �Wv�$��f��{�:s�MJ�6YD��e���s�<-��o.��V\���h�+�L�� ��}m��?T+�kwgR_Qt-�y�����F[Q� ���@DP�:����J�f���Ш�0�,U昚�-4؊�)�z�C\g���u�)t���GO���.C}x����v+�ܱL�g�6b�����.�^v	V��_ӎ�3���}bKb��*�K�(�k�C,x
�8�������%r8w��#���Q��L��\Ξ��?=!��%w;�bpN��� EUZ�%�m��1J�X3墬�:	o*	��k�qW��.}��P�Gm�]��ï��g����3���ю��-ٻ�%�����������M^�։E%�BI�%�|�m���ܢ| 2�z���V��5\�GO�e�C��bK�'��s����;ܚq��F���;��T:�������mY+��A.y���\���Q�qn�3~Q[������[��6M�����9�&A���?��;�e�GTP�(�5�*��$n"ɥ.ѬR݁���o�������R|j2��7D����U�V��>��3����8U��b:D�x�V[���+���P���p��\B=����<�0t'O5�C=Lx���+H�M.<��(/z�����VOW>Y�`Oѱn�QJɩM���ռ��R���=4F_/��!�m�T�s��a�<�/;`���
�m1�Z�j�p�p!qGd�(-����8�##�$���t�M��t��1)$1ӎYn��=e�����"��;]�8*�$��c���F�h0�9l�^��ib+��0�ng�,�g:�P�1���5]jH.P�3�h����*�lr#��Z�-.
� ��Ec%#j����_H���>	��̞z_�CȐL2���p��|AiK�c����L~�����+��5Iƞu���.&�Ǿ��Ģ�a��x ��'�5���=:���D�M���&��Ӆ��oQs�,��2u� ��	�~��{7�Ty��Ø�ѷsjkz�es�u�=�