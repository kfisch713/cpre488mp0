XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g��o��62�G�_�7D;�d���1�U���ko�>u��"��8dߺ�[\�x!E\ٞi
��t���@�]J����������v�����$g�o(�V�7,���'AT�% *U<��yd��*<�{�Zf��pg�M��۵ ��)E�%��C�6�';߲�/�����^���6R-�#r� FJ��T�ݵI[�38)�V�{��jC�ɖ���x��}�����9w��B�ҽw{2��N���)(c�83�S
�H�f��s�4Ƥ�b�/H�&;P)t�Q_�y�4[�א����	��aZ���:�P���:̆������~5�vC��µ�5=�n�������i�;�گ\��$��o��U=���� @jw���S�7����?+�w�92���>�cn�7-*����8��i�����8��>R\
l��1fxI��q�'�)9=Z��ۗJ�;t��"�ʑ%+��ex����XV-�_E�m��O�?��*��}��ʩp���u��߶����|�����2o~�!�La7]@��@����p(�9)x��G>)F5�kM���$m1fI��;�R9<���d��tot�6�V�}�$>/;~�ѯ� �������;(EPV�B�ez��W+B0m�׬��9��2���'ߺ���xf.���H�י���##�v;�OD�f��b2��x/��;JLn�hJk(�[:�jY`;V]M�v<b�ǙmF�ɒ|m(���a�m�L��_9PXlxVHYEB    fa00    2040�+�G��l~��9�pi{B
���LS;���X�װ�a�,U'����������*��E�"E�KW�4|.�R$(�ܷ=�@���Q�)�eV�ƥ�K0�#�:
۾*����u�Qt=��f��2�kJq������c/��@F�H]�]u61G���͡#q-z�Z��f�^R�J� @G���S~�P�H��Oᱏp7��W�C[:��*�?��~�]����� ?uP���~rZ�2qm���/�����6ȯ��4�s�%������C�76��yT��^
�y�'����Q�����!�P������G�( 7ҙ��"u�(�IK��)	u�#7M�p�&� ����f@󳺇b�HgBRN�Q[���l���ܴb�jz���e �?���"�`$J��W���͖�+���k���_��1tb����~R��n�-[������F�q�3v������PrY���2�v�jߔ*��0d�E"M�F�4ؾ�W�o�+=+bP9�0�e��h�B�P�]�v�:��PX����5�g�v�,��}XBK����O�,;����������[�%��P�!!�����������9�ˏ�)��،}$�q�S稻�2��zEO+��k?nP9�z�i8�X�R���	m<���o�@*a˴Q����������� %�y,<1�_��
���Ӟ�?o�Lٌ|�v�'J�,�ـy<*ύ���ANܯ�@��<�Αm�����0/g�>��j���y�=���΀��ǈez����j������;���j�'��?{tJ�X��޳ M�-sp�*�Y�Ѥ
����������Q�΍�Ud�TC����[.cK�i\����>�l;���aJ&��e��V;�B%I�Er4�ikۀ*X8�W���t;�g#
OG?h���HT�<��%(�P��o�a��@@�J*��L �G�5��CO�4WW@L��%[��`�m�5`�YЫ�*���hO�0G���H����N	�1:�]{�;�=ڇ����ԙ�]�B�a(zl�� �ƣ5մۨ8Q!��0sC���}�tY��0�����x��vJҘ�F��r� �\�	q��nx��H�ZFB`;%1s#0?�8怭],2��d�Y+����	9-4�`�nKzɣ?���8Ki&�ʹ�}N���;�-f^�yI��x}�?	��V��g�Ts�-�D��1r�L��'.b�jΚܝ�P(���s�nl�4�Cf�Jk$Z���xV�?_��/��o?\DMę���e�����Vt�-����>�G�L'ۄV���S��j�3���fB�2ˬ�`�{iO>b���]}�fhF�۾+yH7��>�#9��K>(=�6w�E�j�͘�����b>��IrI�q@pG�΃��Pq�s�=. $7stG�u�r�[���tkV^Z��c3W�u����֞�W���XTtܑ�ioA����w�{.��RO�x��%z��2��k���i���x�'�kf�dx-u�g�:Q�7��Ҽi��~���th�?��!L�e}C�e�C�L��� �7�z�/�r��3y��a�+���Dds{�^P���fLA4�xE��0��=� b��c��4��Pּ��3���l��^���mӡ-b��t�2	r���f�d
�<=�3V-��Xٞ��͝G4�qǋ����L��NE�*y��Zo�ovߙ>4�.{�k�xP���-g��n<��ֈ�D��$�X�J���Î0�(w��k�M�a�V���J��+�{Td&�����:u3c�%��9H�8;�Kz. ���Y�`tm=�%S��la���wL��V�%�I�4�:������7_���N=-�C	�w�}�iT�_��m�˲��������sd�y�̏��ٮ����g�m�!�G�X�S5�
~t {wW�2�_�$°�;��}��VP���.���<�dޔ{���P��:�:]Xٸ����?@X���m�`���Ej�E Nn��nλm�`�O��ïe��S�:�Z��nv����U�����x�{�̩�wV�� ���ʳq���d���J.�����C�{�=�M�FV�3��y�:�i ���L\)�l��T檳~.0�F�`g��^wES����"��0���
\~	
/l$Ҡ�K�ߒ�z�M�zF�K�yK�d��ȉ�l���y��l`�E'{%�k?
�ڞ�;WzL�39y�L`L�/T�I�9���$k(9���mc2�����o�&����W$�g0�ׄ?������$�����?UW��V�*����*�O�Y�ז�O����Ն�f��]�7̣�P�c��ni��&mG�!Q��K�s�1��=�hNUY�]U	�r�@`7:��=�J9!4d�4�B\��9���K_���Ph������Z��~Z߰����*��/lv{qc�a����f�w�a�좈�[�t"�����3Kr�?����.T���Q������u:]z1�L���7�ZW^AnA��x�R��	ˁ1E�[s+L� ��V�0��4�IC���Q�*�;Y�X�c�n}�Љ��EJV`�#��u1y�˟]`w���}f{[�*�P6>��Q!�z�g�P` ư)y�=�-����)?i"�h�.*d�|�h.�X-��A�}�����*��4�K�������h�7[#Y���=��F!�93���Yeb+��Jb�G�1?4 �^�ĸ�n98�
��Rns��:ƈ�փ�)�u��+䝋z���n3X�A9�����I�ƨ�{8Xօ��_�
Y�`�����s(e=@�����0�6*����%Ǣ���wr�L���v�$�P��7#�漄��F! ��>h�$�0M�*3$��{��k�d�}.ioFؐ�L�Ӥ� ��
��@�9I};Ny�
<v����3ynҏ�4b.������W�)��$\ �8����s<V�GԤ��Y� �eJ	Qdk�.��v<�̸-g�H⡰4t��9Q>{�x�����S�&�6Pϰ�O�	@��Y�>[��`�T�P�E�%�I��P%8 ���K��`�0,����8�p�~:Rt�_|7&�#����&_����hPYz{ 8�I�����?�[��OQ�c�w��o+�4���
$��REԊ��iBa���� �qEh܂���XY��*+�L�ɁY?�T+O-"m3Gj����O�Pm%�J�t 3V���R��6-Q�5.F��Ȗ����^/XJ�ћLf���Q�kʢ�]��CIR:/@z���lӧ�4QCvV�%� /�!-9��Bk�?8q�^h����a���(�+��`fГ�T� ��2V�T��i騼��W'{TȶS�R��Z^�'\jO��3x�rF��*ݷ)�����M-p'��E��_^�7�9��CY�5�Y�]6��崂%D��]�4/�]@#�D� `�����G��L�`��hz��-�ޝ�R� L��+�d�-���$g�L�/$�F�ayҵ�G��_"�}|��&��xW��0_R�W#���<���~oZ������e%U�Q!��`�m	�+4�;�#�A��9{�fRL��Z��B�%w��o|?���w�Y��Ӵf�CYP���|��:Vz,� 0���-��8d_d������[ݠ��v���Rl����f��W�i��0Qr6�����l%?PZ�$ u����Oy��n(��r=F��l�W�65ʪ��T�#����L�� [gT��t�+v�S�)g�����}�sf0��$���t>��J�,��.%L�����ň�$�W�-e��X�B$lb��)J(���E�zyn��~o�s�C?��g�>��}]����@�~�T���
����t_i����As 0�r�E�q�PS]}���~���V|�VA��� ��*	�K�q��!�Q�[خg�؞�յ�ױ*Xa�|��K[� VU��'�v��3b��S�<��J�8�I��vY��9�����b)��}�k	MM3������,���>�APT�O�ʨ�C&���=�"��SH�=ՑL�y��Hӓ5ȶ�Ƅ���']�,b�#���9X�\�_��P��,��"u�b��2O��[��M�L\@����Y�z�g�<s���e5����f��c����2�Mub�:O�R�gs�1&G�d�+�/ & ����u7u@�E�g���ڢ��ܥǟ�Tc�,��[�{?H����,��3��<t[��b�'}�!E7��^��1c���FN/D����3F?��wT�a>@� {��t�d'�O^cNC�7��#f�{�11V7=5��'T�3K�0�M��6Q4K8�y��l���<[э�V�a51l��ǣE��+v1���FPK��	����0�di�[��K=X��=�J����	�ń���:��@,k���x���}���՘�����q�ն-,�Z ��dCy}�j��Ǔ(�=����O�?)�u;�+��]�5ıy�c�Lȅ8N.��=�П>���z5���SBHd�0¶. L�q��@(H�k��yC�lͺ��k�fl�0@���,8/�ń77� C�.$sM��w��6�:=�[v���P��UE~ˀ�Ձ���;�u�t'C�>n<b���?���	H�h����a���]JR\f�h8;��c��j1�bL��p/��·;�U��Z�|��<.���_�Ɂ���K�A2������ J�zM���Zx}�L�BTʜg�Ӷ}�\Ȉ:���o�ɾ7���%X�Y�Õ��a�2�\��Ǒy��5�FP����W�v�w�w���B��5W@{��f�+
�UC�l|t��'���! �Y��� ��_!?cdX�K�{��+�X��U��f_Q�s������C������pJ%����b���e�Ns�Pϴ:hB�p���]&X�T���v�Ǿ�^�,�-�o��ȭ�_��Vcj�ۜq�,9�.0�W���[��L�A\֘p:!���i��P�N��(�un�<����3c�^S
t�c����&�ø���џ*��Лf��l��� �r�1�O�Q,#+mC�}�];�gk������t`N����"[�7?nu��1}��VҸl��c@˱k@��؟\�!�U�=�f ��5;ca���N)�����%Z�.s�N���I��=&w�@��tպx��2��̭:�Cq8���)�[�Z�^�{ڀ�C�^�33�U��q)�lp�L��As��'!��7�b��|��M�6%�������;Ђ�R*�E�'�S��}� f�*�`-�i�����QA���ە���-"�UY:)�B��ly�)7>��T�C��t/�tV6{���u�qQˮ~J�@�2���i�V9(-#��;�����74�R��7x|�(!8�{�9���b)�2͓�=�2b����X�UA�����{ 2_�A�����i$�P>���ҖX�"���.L=C@�<#��*r�� yJ*kH��ۛ�~$����{�ԊB���M}��$��D��~�968�c��L��.�Z��| ș6�A=�a�(mG���=s���o��"X�E�H}I�H�`��PM]TH�%DU{��烹�U�H���絈zC'��HZT�h�=d����%�#d�V��$Fj
� 'u��xSV`i�A[��&3����7Xߋ��+7ϩ.F�A�}n>N�%91��2�W���#��'�=O�#HM��9�!T] g���(�X�i
k��9E%���^�Kc���BE	*�Cf9Hz.|����X�l�_*��$o�x�n�$�T����������x�� 6���������2t���*t�*�V���=�� �����:4B,���lQ6!�6 ˺=�p���Vɍ��?��<XNj5� �J<�3z�fw��Y����tf�\��CC%!$zz�`+�D}������댯g<�F�ѵ.Og�^s�$ a�YT�+C�E�a5GΗy8�/�pJΉ�F3e9qh��KE73��t�y��ĝT Q�#�@�����8.6�'�]㒛��_����*���EaT3>��P�����-���B�\�nrGޣo.�@N#"S �%hOE�lJ�db��j�0�7��(G3n��H�K4>:A�i��ה��9�BD� "�K�U�%���9�~t�fr Q��}:~��{$l\R��ԡbJ�zuE�LZ��ZJ��|�(p�|^����z�"���Y�8�Q)n����Y�q�bٳZ��4h�ōj_�&�Z���u|���G��&p���1ϩ(h5�~R4��<ZҌ�hw�q�{ �]��e�j)0}��$��ӻ���b<��=�}}1�.,�O�ܾ�6<�w���o�[f-����!�>N�Cf�7��	��}������{5(5��� g��0�+0N��˫p)w�4��#�Щ�
��GYv�VB��!6� ��9�3�ig�	��4�})DzQO_%)�^Q��σ����l+�X�1���T�+�/��	�+]K�w�
��]�9<ݟQ�������F��Gv-�Q��N:��ux�J[`���kw������K��OX�Ү�A�zv|��u�I
*k�es|�O��h��_�XP���L�y'�}���q&�J��0T)��;6���iC�'(i�Dw�4�w�5%�y��vagJn<7&�������A�
�~�g㽀���cNP]q�"l�똋�bp�nɠ��;H>�@`L�P��.l��`�Zވ�XT4���r�!����� 4�Xċ�`2��JOY�H�	�ys��Hl�r����P;�d�St������������	���{�n����i�Yj���:���`GK+ eǲN��z�^�ĬN*�/+V皚�2�se~Mi}M2H������߼�qY������m�آ������$�	Z�Tb�>��&��?$�NY�����O��_�rF�Յ�!�ɭ?9��f�X��b�О�0��Y^��ή�&�J�#�~F/�"W�����`�ƀ���F7�(`�͐s��� �?����e�>�4K�(�:V�rN�A�oԪ.����.�@��p�H�u����M��%D1�pn�w�	�O<�����E�S���׏�p�_���y8G��a[����f��$+��X� �%+Ԃ-*�`m��/����Ú��(`
 �N
M�5���A��%Fq� ��gAZ�+y*�E	�hu&�\py��ǝ֗=��
���[6`��)�D���6�̥�mgJ`V��:�u�K��,(�	�?tdF�6��K��3�G%%�]/v�.I��p���6h�UO[F5���H�Ӌ`�Ĥ(�55vW�N�4�p�£�MR��;�S�\��wN#��s�e��m	���P �@$��uG��=q2�6!�xh*jS��-��
n��TǜQ��/Vl�d��>�Դ�����:�i�9At�Fy�XV��5ld�\7�pXU�٫�8{�M��ΙN�C{V$&:щ��m=`���ߘ׺�h�ȼ�������|H��_d%�����r�%����8�%��8����Dv~OEu;q/l;���j��#LkTbƲ������U{,O���e�CEc��1<"�X�ǜec�Ӳ �at�N	�ŀ��T���Ǌ�u�.}~Rʊr��2s�.^�"G+�p���.�t�	���lS����`9��i1�ͭT^*8�<���?����IV�}����'�Бґ���:P��U��\0j�� �J���D�	��[,z���)�@��ΰT�����\l�恰��`�^bՌ�Na�0��K��;�Gƅ��&َ�F�"��4}.��7�B��;�����_��p|!�R�HY��WVe3�&`	T��P0
�g�p8��d��R}�&k�%�C�:��%���B������e�0����)@a�J\YlHu���~�q��{� ��e�i6���؏�_ͧ��N�6����|���/j!���,�س�:�q��0�O�}V��9NCй�O����8*���,=Y�R�'ʡ,ǒ\��Yj|o�DJ�{,�z�S^��ݚ�5^�n5�Yl�`Q�ޡI��E���w�-8볰o�NhS�A��g%�;ɘ`�ǿ4�
�Q�����O/��F��N�.>��P�J��s $��P���r����M�'��^4��|("�qM�fXlxVHYEB    4f62     b50🻡����Z35ܽ��Z�&���)**Tܯp�P�&4�}w <�֥�Ym�CuE>N)��.L�#�I��t�v���#��r��3�d�(a��L���,^ţ�+�\뻳�aMł1R����f�-�(u�	�}�X�� %���wLg���2��� ���E[�j=8 ��*��\ ��2e��>��4��=P�Uw^=lP��븷0��m��{p+?�aKl3��w�Ŷ���I�bd�6�j���a#��b����ٗVܤ�&�X��a1F򁺾&Qc8$����y(e���_X�$qԣi�ﳛ'RI�Z��Q�b.�}u��EL|�ڰ�^�l
+��BA���&v& �w7�V~J��}$�f���Vo�Ht�-q�=��v j&�sMT�hDT�vX�B&��9������%f}��wl��3��eP��:͓�	$eUcS���w�~ WOO�ꬭb7�ve�e �`;TgX s9f�9�m1i M���Gt�.Cz���q�$:��-�q�ｉtx��<�J���fg��t�L�$��O㘇&�=� c#A�F��
��x���d�ě���{����O6'q{�&����C��~���W�3������)U29"P�/��kZ�x��L�f_=L��X�:�ձ�>�y�Iq��	0ߤ���L�.>��X�;��v��� R�뿮��!4Akio�~�e`�&��$K�i"}�&H��55�f4Z�+�(F?���I������(/Ӌn��k��npw��_�t���zz��D/��;%����_]\]�h
�P�G��l�X^C�J�7����n�]�t�+�R�Ő��n)AlX1{O��yOEP���p�N����1e막� �kb��@Avm��\�{�O����ʔ�|�=zƧ͜����CCH[�v�$�gx�։H?
�N�u?�����(j�?ܐF~@S'�fr�ިHH�Xde�UX��g�Fd�Wk����?�5���)Mb8	��F�ت��<1���`GF5{���fW� A;�m��-BQ���mV�e1�|��?��x_�{����r��Qa�Ay&r�l}�4�E��x��R�����+?�S���H��0��{HN�e��P���\���[���?��>e�Ɨo��mjb��®�y�զ�AKo��	{��0�mw�F��cJ�K7� ��������3�eC�� |:!�IY�--.iݣ?#�`W��(\	攟I�/y�|�~���Ϙ ���8�Z ��	2��E��p*�K��@�Ih�]���lG�����9�>GD�j<�k>�՝ga��o0�jKv�A:����Dw~��J,؊���HC?g���mk��ڿ�!7�T�~BƠ���,�b_Ⴗ�b�f��_ع���B~
�g���A��]T;؀�{̳��{96�W�����_,��а�b19�����<���%$���/���h�CK�v�t��P�cg�Y{��O���<�<C�nV�(��r�FI�2�9GRDi���˳�z����F�/�l����,��$.$�P���}��� /��`�_m�z:���}1Nv�V�z�� u�R���mz[K�d��Ey� ��~7��Û�#�7��दS*�r�5a� �7Xm��Puu�3�h�gL����}AN�)�ʏ^�9]����5Ћ�x��ʚ`5�;�)!��1H���	k���M�r�j&�yE�&c���D��\��Y��M��� �hz��&GQ	P|�ۍ3�wENQR�L�#{A/%Z�����{k%l��\H�3!01+.��5��7t��������UVd~7��X�/%k*���Ӹ�ԙ�N��$Q����Ö)�Hg8h �;�\j�FJ�w�W��ed��`��k�����h�-P����. (,��"1�_N�x�ˎ�L_�;Ǌ���N���[��g�:z���1�܎��}i������5g���?U����/�`��!]`���5��\�S^�q���F�K%������(�S�)^=)��26�����2�;r%�k��{}�˝l��=�W���3���B������)��������|G��	�c����q�Qڬ	��bJ���� ��,85fI?�M.ـŔY�(�!줽�<��A,[m����܍��6�͚j}�~��y)�khW,f����N�w<�5�7p=q�O���;�KU��2��
>	{H�;y�b1q�ء�O[�Zn6�W���լ�|G���9�	�1����V>t2��r��/<�Bo-�33D����JkHSb�{��Tȋ�d��������:/�Yj���R�r�*�#���_��WMB� ���f��'⺷�L�\B����=�Y�:><漅3�Du��P�Ĥm�E�:n�/Mr0T����*y����v�+^zs&k�g��WY��T ݓU�~�'��(��^@��&��=�5��oX�r��l�<���|w�bi��R�(A\/�W&G����h��l��M�J>{I��_�\j\�%`)5��/N�ndv9G��K�e��
���;���8g!�ed1I8��eƏۣ�6�C�`+lB���nL�6P�:�~#XȱE��Z �ͫ:b���׭��\�.��K�	�w7�v�ۚ�?��MV�z����\�%�����Ssٿ�-��}ú�4�Q�����a�� 6$��.an�}��ịiR��#zf��W'�B�XR&m���}0�֕�ѹ�2�5�
��������͛
�XHxD{�c����Y|�^q�W�Y`��Iܲ�L9m��x�@���V���p�)���8�����Z���й���̷@��e��:e�T$[Q�ܵ�*����� ÅA�8��
[���hY�ck��