XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8��z�v5��������C��~�*�^?19,��I�X�bk�7�
C6���2Я�I|���2��l�v���uDω�#�R/.���@�8�u��:pW.]��xM��*a���D��Vm��a���P�z����y~�݈Vfid]
�2(��_^�v'.X�Ї1��2�T&p#��D��Ի���?�=󤏲�ȼd&��:��Q�^���Ѻ���e��u媿j����݀�3����F�*Z���:���_�V3G�Ñ�(P�P����Z@
��Α��qZԉE��</r7��=���~��^���� Zy��RɃ~6�<fH�]�kUr% � f$�#g��I�Ue>��r�FI��/�`4� �B"��;M��F�6��=��ꄧ����ǈ�_��BI�˄A�	d!:2�ּW�м (Y@t���6�Yܠ�Z[T��YQX�Ƭ�c�Y��y�b%�D�?<7?R�X}B��^m�Y��f�lR�iTY�$��vM!Dh�n�i� �P��L�64����Y��D�W���l�:���m����k��9+��I��H���Y���!�ό'-�,@	���g�iO�bŹ3%���\$����9������^�#Y��q�����h{u�c+ĭ`C���L�kDD�}��!Tc�f��LVf��mM�'�Ȟ���K��㕹�U��xl��y��u#t�i��$�|�YDض���/ro���]T��`���°���Fi�@,)����9���*<�XlxVHYEB    95d3    18d0�����{ AkZ�:���7=��Nw P�%&2s,��p[k"V�$ߜP{WPtp����q��e��,�>4��x��Gd�p���� WH��OJ�2�x��o^Q���!��J�?�Ȗ�2�6���c�E�+~����$@\������	����|Vk���)K����U6v�a��u�QO1�.�嘛�,GR��p_�l*5����X�:��> m
3�=�'�¬�?7� ,8T6l9���t��j��>F�QkA1����(�ndVK.�X�U�>�@Ő嘧8KQ���4G�_���k����0R=�hP���e�=QB_�tl��P���6?]X<A��i}�뙣@��'�i�/��	o%�'�OmxzLx��M��	�����3�
L��!����vD�Y�K��"�&ErXL��"BKK:DP%�J�h�L��I�<P�Y>�v�2��L�O��$�^	������)+����j��.O�m	��Nn���|ѯ�X�� %8�`������ԉ޽��w���Qx�E�s���GF��v�9\���_t��D'(e�?4t�	��Ð���߲f�a���x<���� s)�Elq,��ߛ��������Ru��*�..���sұT��k�¿(7�s���ͨc{��M͢��	a��+*��BH�v�Kre�%�dt��O��2$�&%'4�� �OusbTÀ�-��O���-8���0�fT���,c�CW�O�k!��i��^z�W)I��\�\�@���4�����7��WS@�܉���u.
��~_'����^	��"�7�7�Kʽ�1���}P���9Y���Dq?_y������o�D��>^���L����T0�<hP'ȇa�G?��Sȟ��a�?�(�	����P�wK��v?GBM�����#�V����0�>P�A��q�@O���%Z9§	����L��<H{�e�YX&h:5b-�~�#��UcAs*g����&_rdP��/�.��*��\�����r�i �\HvpN�D{i�jv���D�V�Ѩv��%�v�/��Av�>8g�G�
�k���cw\�!���X{��;�n�Y������JjPoS����޸ �Z���UPŷ'��V8�l�FX��@�QF�ʎ_���#+*jET`�n�hx�+���������a��EN��{��aw�GzI}�:K*�W��^q�<m���N"KR���Nۿґ��Z�2���w�\�u�*��Ю��=�S�]�I�B�h� T��Q�Ξ^�7鄂��xKٻ�B��ɱ2�.7h�Z���
�rM;U���`�i�fw>���������S~l|�i`�1}CV�Ĵb���Ü��
F4�����:�F/� 1��'�@�������Q��Ah�YE.�+�)�j	�C�x��,�� �Q�E���N>�3��x�E����;���i���0� P�B�o1����#58Tk�|���ߏޅ)���q�\څI10�1�9
�C����rJ�>-��㕈#�hY�F{v�
����������@#�҉d�4]����=�5��8Ƴ���NP�(��k��|�C�2�ik�>Dk&�k�:RtS-0:�����1�\�.3��фY h�(�]$��s����cs�|!!��|ꅃ`%���|eU�)/I�p\�����O���s��饒�v�����M��qtK�P;83�8�8�[/��i�D۶d�3��{{"fvL���ib�V�9g>�H�b�ta߂������ƑNu��p������'�!q�o�?�j�lҮ���aV�^�x���(��FVN(��&�>��+��=�J��:��v@��#cg�o9S%"s�s2ݩD�0�pO���|E��c��K�*N��3α�6NV�B��u�������3�*���D��
�+��g���]��>�y:��j4�Y��	*S���Ag���C!<:��,C	R����-�,=k���K��fDR ������ܜ�̐�@-h�k�=^	WU��*"3�/W]��:��e��m^��o����t�b"�&�=M ����`�#*0���,����)D{��l%��9�$>Q��.�X�&�1���������EZ��h\ӊ��LA�5R�q#�ȧī�A��6o�]��X�"Ϭ��֟�k3� A�
�]F0��D�ti�G�!މ��_zB����j����j�)��< �pP:t�K�GO+�B)C)z���\�D�-Y=��dpE��2����VGJ%U��N���T,S��$��yNG/2W��� �>�~��b����mZ� �L����� ˖eU�h��ޯ����7v��f�6�����iW*�$��ɹ�cs�k�m\�-h�C*
w�0�7���Zm�jx���A�x~Fq��G��R����	ؐ(�h�]7���8�(�'��U�_�� ��J�~�@��D0ԕu�Z�=�#���.�:͚~���@g:nLGOH�op-��~��/*'(��v����p�M ����"���.bpv����.��%/��8ʂ��tI�����p�W�jj�	�R1/ʶ�U�H�|34���F@�8���'��{킧.�X�imT�7�ȍvZ���Hilv��8��8���/���X��$�"\E60]������Z���ҹ*�j럿�i��^~���k��B�5�ř���b�j���)|�/n���n1д�FM4�O����~f*�^uXȘ�rE����w@JwXzW,ǎ\�J�Q��.���I#e�ɐd����8������3���	^��>�ˇ̈���/�hv)PLZZ�F��"Gr�=�7e(ea}�}fh	cYh��}S6��k�8�ve��}���z�h�V��sz�~�GG��iZ������2�7%h���b[o40HsH@�	��/梴$�?�J�㶬�gEi4,Lꗆ�h#2����C��(�R�mDQH�&ʓ�>���a�H���]�_�e���J�B3�+MʆYdc� �6��<)�g��`��»�d%}���^��s>m�Qſ=�)�̸����j�lABC�oH,��2Gf����"S!ppU�5=�����Ng�]���?���|����$Ph�e]L<*lo��"A��g&.����zh1^ZIL��Z�/��=ŕ�hL쉓��vts������E�2��6���i�^�8� ��z�O:J8u�#�C����u(�#�U�TM��9��f5��P$�G�i�ѭ(�Fv��)�Znr2���3�^�� �)	��I��O|%���W��&|�aRh?0�`NV ��w�k�1�۾.����I{-�܋��Q|�L��MN�h�l���Kt�T��ՌiY��_�p�ͭ��+�z����w1F����@���tN�c�/)�w7�2�ԓ!-
�/�>/����~�s�r�e�z�J`I@G��d�R�Q� T�S�G����~Xf4�3�4�Wl�(t�p�����h�1�L��P����"f��<��e%ݳ#�O��*RndG/6T�e 7�7(�/����+�$�T�YF}�a���i
�^��3��S�f�� #ϒ��h�f�f%	^#��:���#h�WΏ
��z<;�~���6��]2z�U�l���8� �ېu�AS��s=��1�$hD���i#�a�b�J���@�F��>"�E���8[��u�����~6��baJa��㏒�b�c�8;��z��(p�^��l�&-տ��O3���"�]�K�U���k?�g�8|���|��ȫ�_��Y�R�o��
�L/!�ON�Ru��:�\�!�.k9�
�PV�="U�@�h���i/SY��\�M�G������?p:_��.�eg�雭L��o1�)������$��!4r}��SWW~n"i.�t�*�1�$������!�, �`~Bϭ�᩼R��l��.A�k�]0�5+�YQ^_���u��|u�t�R	�B�����z������a���Z���d@�d�_�h�T� `�/#��[ZF�2:���+C��@�8��-�`����e��?�L9{B���g:k3�p���%V�0sa�����HV�F%n�\��ΑM�M��bF�W�lN���4��T	N��'s���
���6DI(nH0�X�����o�th
���P��5���نkp�<�x�u9Ѯw�ޖffl�~��;��Gt���!�'��U�Bd���@�D�2��=�8�nm��CȑaϷ܀�W�F�2S�^�+A���7���Uqw�{1n����=z>�b����ݮ�X�gy�kI=u��S�7��q��w;D�H���*�3{F=���-_�a�D��U�ř�R�[�X튞��}K��<��N�ųt*�z(�P4����6cx��^:��ѢZ��\� �AУ9G�1����ϪQ�Q{՜@�V��m��͋�;��^+�i����UM+Qa��-k�'��v7�B�T_�t���Po�Kd�L�5K$�
��`�4^�(:���1�����('�a��_ީ�Qx�K�ԪXOkZ��Vi���t�2W��$�B=�����P�*��<6.\߼�i�AB\W��h��5�������=E�"}��vx`�����4�`�W�s�n���w��;�r=>g''�Y��&�&/���vNGX�u��Ҍ�L"`1�-�!a�0�>��|:(y~�#�휝�p�~m��Z��/b�\e��7v�,JZ�_���Y�FZv �hR@4��(��J��T���Jt}�@�����[��Z�B��k�}�C������R�}�B���C�tQ W�I(�@f��0���p
���>�|�]cJ_&�Q�6HW���S"��<�ko1t���}ΗL������S4��6�:�?�i=i5�j�G$��p�5� `[M`貭P�k�#��t�<G,�j��ހ!+���eQ����ER��7ꦟ�#��Z���=�,�,���s��~��͛����hʋP�=��k����sV��",��@�.O��mM�������Ĭ���������vq���@�$u����!"����� �fS��(�釙HZF7I�����<0�޺V�5�g��J6<gd��d�l�L����&�~��|p���.�^`N�=��������!k���CH���3BF�A��$.ch�.�S¡�����Q�����-�)׹�΅>"q/7Mjfu_+��� ]���@k1��t��c놤FeJ�ݳ��l�2·�~NU=�S;��brfq�A��@�V�B�� H�&�6���vt(B�n���hem	��V:�}Ҽ�#�~a�>��;��F��$�&Fd��H�!V`s��'����+P�+�8�`rfs��:4G�%dԋ~';SJ����P\`� ��̢�[���J�|3��F�?$�˕@MN�Hp1���`x��1�/����k���ȃ;�`����P�訆jk��|zc�E
�ϵ� �](�����]�I�{8�d�X0�D"���t^�P�����;�r��-�m�� �e&Oo)ȿv1GAA�5�ރ ���������1:�Y�L4��n��䥭����zxa�j���Q���f��}�Of�>�;��y�9:Ğ�����JBbS�~DsX�0Χ��D�a��%zۢ�)�j�;���j�c������Zs��;rT7��Մ3I������z1�NgWh�̨�Dv̼���D��"���ZEh�YH�(�[����O]-/�_�D�p��8���b#��xGNȹ;��*���f��IAgy���ܰfZ��p'�Y�U����-.�p��H9K+�.�:Е����&����R+V���j饯�P�P��D�������uQ��YO�N{��arēԣ�r�d���q���F������@ԇ���%"係���2�,���q52�ޭ�,�oCU�6�������De<x�&������6��!�K��>-^�N@��Ěyw����B��_�}d�9�h� ���b�-��!7�R�(�/R�*+z�TN/��YN��O�8D2�]��	�a�|iK�L#A�BÂ��oҒ2�~F�t��\��P�m�`��!�+a������
�	��R�v��	\yvS���.�	��	��/cl^p���%̰��"������/Gՙ�,��d��LIv�yE���`�h���<�hƮH���w7���	�%x������/��&�����������#j���}t+��$}Ƴڨ��Z�V��� �1\��!bI