XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��a?"�%�S���4�8S�u��ض'�}Ϥ���:� �O���0��sD���PSU�L3�re��o�U�[ �po/Ǟ�Ғ��~����-�#�L6'��{��a������S[O����u:5�����%�żNɄs�������o~����#Q����;�#6��VH�W)�iuA9V%3��S����\��E�a�5C�IJ48����!�HAG� <� Vϗ�� �<iډt6s����5�Ü��}�}Gp��$	�xZ���QN��G�Z%�����P�_3�s�6����V��-|������M�I�K4�A-gw_�E��
��P�5P(���ymCB�����:%
�Vޮ/�Lv�,c� <Oz�c��o�`Y"�Yl4 �p�_�z�T�d�$��o��{'�I���)XJ�������6�jP��aU����;�O"�T�P�pL&����빴���y����L<R�b2?�$:��`"-�E;�r^��2�l��&-��I,�[�#��d�����폚^zt���{�O�]���,}�5I� >b�lk����`���:O?�å���X�K��'i�ƈ2hw��<��[�:ڊs{7��3�{Y`��u�q��*�����&���G���D��N��F��k��io.D)�2|oxS���[nT�^���F��3+�h,����D�J���Oae;����X?o	YRb9%����ʪZ�
-B�����L��c?t�����XlxVHYEB    a037    1fe0��^���y�Յ4�/�`�%�.2}�c������E0��J�%E���r_��퓿�5gx`H�(դ��{�4�9X�ˏ1n�Օ%�r�:�*�T���S)d�nB���]Ld���b
���L��������M��荫�k��u��s�E���T��Ӌ}�`q���m�����kA��KKa�,�I��E�Tv��	؅��6S!��z��v����F��������"q'I�'�Āw�� ��s'iE���`'a��L�n�`����I�yE��٩�TV��=�D��2�<�!�kZ<~,:��m�I�u���W!���zW����*���*kU;%/Dd&WqiAU_=�U��S���e�-�w^e2��vx��pN����^��Y���c�����2�L
Oȕ�^�G�X���#j�gLS��1�Q��)���E�
ฌ�"��"�m�G�X���T���>ye��o_�Ud�x[�!���Eș�k�p�X�gJ�f9���2��v>D�#��N�y��N��P4KG��Bdo=t"7��W����2'h�㑓����"���7Nc�r}�
3]%����elj��j����ŧ$�M�K�v<��X�Q&��G4����N��d�p{.Q�;,I������=����v�S~�]e�Iot6�a��ite�e�TCQ���Ȩ~��xc���ˑx-m��s{�Nj "
���u�b���S����م�8���2�WS-s.�~�`���hf�Ғ���u�Kj����n���h����I�zD'��ck�+h+��kcrA�xO�>{��ud;5)`�gY���N +��N�r߹[��5R��<~�xcS
���F���!�N��i��y2�qu,kx/Ǯ���z�S���F1|��p[�xk{g��s:V?���)��uOy9�m�R��̌~6
�S�̅�>�fh��kO�j�D3�����^�����vݢ>E\ vV�	o�A"����&�t�-�5��9fi�Ը|]E� DY��o��(�E0wފ�|:�!|��0�AI�l7:&�,]S�W�tC�D1� �"���Ѽ�M�h�=�`�������!�V^�9�({��q�TD0�e	�qˡ&[�Sߴ
`���>\�7]̀����n���_�
zLR�Z��G���u���0���`��������ތ�Z����{���y��zʯ�8�i}�j��eg,u��A�aɽ��~Q'�3�	�[�xn��߮���>���n�b,˔I��=�0�6;��7��z^ZB�1����	~� ��|���$C-�*��`,��P�7ب��ly#9�M?�-g�vط�װ�Z����_8�٦�-��"����mωA���Q�>�%�m X��&�]Y�P�'��5Cx��\��=�},�_�H���m9��wj7_��n�E��s��$��8OX9��z�%6M/���D��l@n���_'�ݮ+�,�<`0�������y	��z��;��k���X�N����T��H��v��vx���]�Z;��K3�<�kX7��w7?MAR%�l�m�P/���ː�"��w�ۀ�`�ypʣ3�r$�v�� �XG����`��v���N�$�dR{�?� �C�,s�����^*=+H++���W�%UL!y�S��3hp�����#cO*��r����łq�k�P�qr�!��7��ۋ�b\��J"�����U�G�;w�A��������{ׁ"��������N� ���Uk>ͣE�߉ ����+���+�4�h�ⓐ`��:��!#@�&��!,�&*0w�Ye�Fώ1EN˫� �%t����p��L����-Y�G�^�LO�L�b��:��J���0��DQ��NR`��FO_)�N��(!��>�'}�i'8��<���fN� �]5��wo�9g��w9��3�������N{�[�>��.�eН_��S���v|��d430�����  �eX:Z?���
7�e��u�|�K#FV���Ⓓ�Ƿ�ȥu"\�	�e߂<ܠ_@�D/ߐ|�)������꿁!A[Kх Y�����c��|���2ڀ�s�dH,/N/�CtL�Je�S\j\�g�q0�U�(G�&����L��2���1�B��{򌅉6�F�_�E��٫*X����=%�*ZX�y��q �,�j���������H;�y���M�y~tk6k��1������e2�`�X�zv�D��$��^c��@s3�8<��:���&�q\�qR�D��^Lp�]����V�?�����N�EV�_؛ȶ���E�%w�y;�<��/\���[�|W��?|:>���j�����r¼N=�Y�7���06��9?�yB�;C�dX����ʊRԍ����"d�T�Mv )z��D��ڂX�������� ���������!q_�y��CAo��[jɚ��KΛ��Ly���jH٥����r����XV��P�iQ'p&�NZ�}��:Lw�0ǲ��
_Imy8~S���a[���\<޾Q��O(8o�󇺵=`Wu`lQ7�ش�&�'���m�J:T`��l�[�B[��}��	n2L���ْn�p���˂�t����s��G��ֶ9�e&5b���ˎ�׮��w�M��fv���܋shc�^%�$M���Bs9�������D�"Ę=@��	��A�?��E�I�r�+���r�Ȁ˴����~�@�i,��tXL��W���qj{R5t���'̧�	j�s���3��HH���Y(He��K�8j�ʜ9��t���X3OE�Y~79� ���k�n�bk#�M�W��So�r̈�׫5J�?����{_[u���y�q����?̾ˑ_�<����S]������=��X��Ya�qR���Xt�8P~̜ti�2�gpQQ+>��V�ߤ�e�u�)���+"�CO�Do��2t��*	�����:@l;�Βw���L�h���:T�����w�*�Hg��3⽀2�Sp`�wI�sF����lsf�/�������Q�5v#v�7C:�.s�����
uхF�*��Sl�Z�C�c0�\�O�a�
p2-`��Yс�kB�A���k ��įڲ���E�*�����k������C*\�9[2�vם�ռ�5Ȓ�6�ѡ�N]7[)N�̨��d��~
�m��U��]�cB�,�ݒ������t�D���\�\��-ҹ6 K���2/R�?�6G~JT�+��+�Tr~u������u�0���26���r�o����6�(�<����)hD/��_Dz]��U������4��壥]��B���5��+>Q*� �鞨�ڎ��TR_�u�dnzF��(o����
�6"�#�����!�P[Aڪ���`�f@���9s�*���j%��Ϟ_:F�[�̦��ϤP��u�f�5�Y'@���֔�\eBO�"> ��`� t�z��}��x��3bs��0ٝ���p}흅Q�֙�G�|�����L��rq���aN��1���W=��-!��mnDiM�Wk?�u8�u�~=�H@�ׇۊŚ���U�:���qno�>�"<�-x��z�o�O��^�F]Y8A��!�n������r�3��'P�V��{F�ƌZ"�����a�q�Q�Ż�<���ź�R������$̘n.�LN���K}3ȯ"#؇�Ӛۋ��R���x��e��@�z�Ì�'z��U[=Q_��~/WB{�f��[�?Gv�R��ܦ+��IM���h���ɨ\�;�'|�N����:./nJ��)bg�Y>)�M"�H�f��Y'F����U�m��me���Q:�����RjfQF�-/��1\c���3�3����E�� ���T�{��v��[Oh�`�X�-v���Y,��W��wq���O�hiJ��~��Ҕ�,���%��pUkz�C�O-�@; W�."OORȑ��a���W8��&ռ��/z��1��\�o`r �.d���n _-%��<v�TLʏEmM\��9��.��� �^yn+0,�o�Y�%�w�T�X�j7��p�P2V�]%l��M���cl!<CV(�	�C�QO|���^���&�m�n��SL��̒G��ZR�[��r����0���X��7v���]�ĠH7\��V��
�~�1Q����� Ä��Ϣ{�R���yZEt��O{�`)��ٳ��� 7��o{�z�r)"��fA+��юJ;��nF�Si� �\?�9請-�N۾ɵ�@�.�z�������$���[>Rj/"�E^�U9堽1!w��E�S�Y��EPbB[Ќ��dK �뗝qQ�=�
�P��R{j��|�g+^ҁ���@�����F�X��J~�&ZQm�"�0�u�m�ԩꃂ�]OƳ��2����?	U#���-v젹��W�����A�"���h�I���~�ʯTԄPӖ?�.K�g!dR�!������ߙ�O@$=A-��Mύl���_�[iI����<�L���Kg���}T��Q�����cz
�)�.�
���6Y�`1z~%)f�2��cnA{s$�������b�`�FY:=�0�� ĬNU���ӝ���n8�(G��=a��<;p�>��zc�Y#����-y�Zf^�v��y`�V>~ϥL���K�e&��@s�
�%�2{�J�9�)��mQű�q�b�i.��Uw_������গ�-'`�a���i��f����2��>�B��5�k6��8�AG�E�c�~�47��H_�ȓ���\1q�{�ĉ&�(���(r��aKT��0֭
��b���Ρ��/x�|
p�י�_�nպ��{m[>zK� "��f����C2�)��y�^$;|���F��zU�	��|3��t��,D�21mAT�=5r�[�_2��z��tIn���e�P�^��ɟ�MJ��^Hhfh~������rH^��k(��*Hf�2ل�JT���
�+�xɽ�I��ơ_N�d�	�j"	��M��IJ>_TH?^�$��q�1���}<-�|�<�u]�"P5r�@��Yִ7�	?"{q�od��`�3�,�~�)�SF��s�|�4�	W5�DZ:=<re��
�ܡ�2A!�s�q�\>%�vLG�U�+��=�9=:z��P�4�Ls����)[����ʖ}&U�E�lð�7���_s�#��,�_�x�ݬ�jh�?�¤큊3TbD}��8�X����}����;�(d
�M�#c�4�8m����]ը�]ܻWI���1��D�������\�=*��d�)YNM��[�? ��R�!ʝ�9�ͅ�1h�߅_^�S�(0�1�я�6��K��1="�A�l陝�kgm��2�ߞ,�[ih�1�˞˓����&z"~bi���hڢ��	x�:ht�Ls��,m�f�V�~q�5轖`�T<���;�$����٣/���dN^l�J�V�u�:�詆4�k+a1��,.���B��FnK�a� ��\4y
�ʊ=�+���GbR�����:4ռ�+0�a�q?7��=ψ��lz � �k�|�/'li��BMF��Q6��׼`�����՞�9R����`2f̷jɚ��^6�3v^�o>�}�ɽ������������v����]eU�w����A���m���;���K�D�9�}-*M�t��Tz���i�����nz.���y�C 'H��c� `cE�gA�
��~?r{�+�v&IW��Lo� GA�0�N�J��p���s�s,k�{]�x���*��$�Q��G��%����V[�����rB�c	�V�3¿B�f*yO�[�\���C᭸�H���i��h?f�B��u=�;� e/�o�W/P�k�����-G~���΄��]���>��(�qg/t3|L�������h�L'lt5ߟ�}�H�uR�n*�8�+��	"���� ?S��#MS��4��d��{ �)-P!�
	�u܂�߬���с�5�ѽ�(G:jD4#ϗ���zR��'ռ�4sG73oB������Y�m�L�f����acfp��ksfŴ��3Z	*U~�wRa?,��	.n��%�^�Ř���ޏu<R�[>�}�_���ϑ��s�q����*�E� ui����d�k��Mt/��H�z�x�k�[�+�6��;��~�8��#ݮ~j�%"����f�!��N%٥�F�H6�w�ih��K��ww˙��I7���@uJ�r��r�9ɍ�z!us�G���Ի���tU��G��	���j����vp��:��G��*���� /��.'�&��Q�(�n^�y32?>�B���<B>G�M�"o�3�E�I��A���B{���j�	;X���s�8�ϥ�QT���>l�!��0B`�ŵ ��ܤ�[�G�7�I����Pݐ[�U����o��g"�¯�܎d';-6�9�0 �R��BN����f9��W�5U���}�<�P�N���]z|?�B+�#>w����ꐜ���4M?f@C���h�ֱ�IIY����OR���(&J�����\ {<��������'`&k0�	�$�8&!G ���6�ˇ�'Ô		���ѳ�ȋB�9"��s���p�T�cu�Q�m����Șg���j�$^��r�t�J�#P��zy�?��5V*5���Pq8��+A�Da���g�.9 b���@��+,���S9��W��c}ejyQ�m�J �P�8E����K���,�KdE�#�G	`va���ZQXP�\�;n�E�t�"��bo#N�ү	b�6�#�3E�v��O	e�nAD{�b5�.g�_��z������ j\�0�7m@s�^QWh�0����^9�~H�_N�C�z��@c�}�Y4yohy�84`���\��.�K�Zg�WA"�����TQf���9}�~�/BC�H��T6������"A�����C�`�K/r
�U[6��gء"{a{r
~����nC
��n}s�Vm�g���M짿<ږ�ac�F
���;F����#�Ĩ���� h���p������޶��U� ����	�UH�l��tXs^�DVE�2?�7ğӎ� ��cn�S+�*@� �^��8�8*�"Sw�u�
���@GeA�O�e�O��^ft�V���q���X��ளD�&b�I��	��_,��#��B}TJ��4�h�a�A�NJ��8v�@aI�r�[���<�Xm���q��Vіf82��S��w��h[�b3���K�V!�/A���@-F�69ӳ��|������Y��,�K�Q�k}�Kp����8���gԏc��:5�����n�r��RJ��ʂji�(թ	�R��������6��"�r��Dׄ�az-�oduQ�s��E�=�G������iֶ�,Z�|���V͏!c��T�P ���8HD��FW(=(Wh��� dG�f�A�&c8�qM�/5]��^g�|�pף�(���|����W�x��H��w�RW��\Ƒ����S��|���-��?������o�I ݂�8"�r���"��/1<H:��~�r��J��}?�5d���:`���E�L�QN�;Š�R���9(��p�~���Eϻ>{���o.��f'H�Q15O�AS�zL����a�7�v�:�8����>����x)��H�w�P�S��Eˀ5���QNR�&v��.z�`옿���h)�s/?�mS�������32��E��4�j�0�i?_�"�~10"���_�3Ö/�L�=�Te�ؠz~�<d��:�\U����0�H4%8�Gj����-�`��,}5�Q��el�����:5��2�3R�nJ�U����9�K�� �@/S��q(i!����1M��Gsd�|j�ևL����-#s�3����9���9������w�B/�7N�^�Ľ9p�p��5
���ԅƍ�r.��3snCy�;K��i=����@��h�s���l�l��t���s���=~T
qg��nXMV'��"�>=�'����$������K��p��\"a#څ��4ύk�u���ڡy���j�׫sy��cE_���	�о��͌��{D�&g$F�C���&�