XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���~J<)�X�H��S!���Z��V9CI��5c�8pb�+�3]��gY!x�ז���g�H����2��Y����>��݋ ť98���ya�pP���ɦL�����!��ڒT�FΑz�D�n���͜��ݚ/v�"
�y�=FS9:��'�zq/�rz��`�d� �{�����=A�{�Z^P~6��r�B�_������l��U��/dM�o�fX��.E���*RF���Xb/nT���"���C�c�1��m�"�����l�Hf �4��9�,yx҅���UKeh(�-y��<Cti�Aڻr-GTc��!���s����
����u �=#�`f���C*��<M���˱	5�>��^��\~�n0|���H�`K����aV�F�-�����l�M�q�3�<@��KH�C�P�:�Y
!��ۉg�j�+��O�H4|1����3>n�TL.����6�q#E�]���� }�%N��7]%��#��k�:m��V��ÎY��dZ�",Ge�����p�x����"A|8G��9-֦k�:�cA�G�ob�����j^&P�;˒��d���_���]����o���[�n��Q��=jq��iM��&Z-�ʊ�d>>�� ��E����V�� Ӹ���.��������_h��I���Wt������K||BE3��~*���cԋ� c�,�ڈ�b��s�%�L	� \��-_���MU`�yJPg�E�N�*/�=
sr٘>�&����J�'j�_�2ԩXlxVHYEB    42ae    1110x����z9{��إjU|�����l���,Ax��l����i���}2y��4�*���Җ�n����֑m�W�pYm�"���ӻ��9��)aK����f}{��1IG�i�
��rls��
u;V�������p�Ξ����|T>��"uwiL>
�����:��U��!���0v���/��ܟ����Q��-�E����|I��ᓻ���%�c�q{����P�ο��ꕈ���u�����J�q.h@ܾ�q����Y׍[���*��p��p�p���8;�?X&<ǹ®��ק�+�ty��;�C�L��O���$*󲠝�����r=��n7��?P��%�mR ]p*��^���˲�8#�c��068��8�a�;X�Y*��!u�����ȑ�xT,|�hOnQ�N�/1�:�%�Uu�'ӽ2�lT�:����߼x<q��Qu�~w�uѾ�*���9�Z�ŵ}�����
�?�D�
�|.WI�t���^_�-�J�c>�/Z��yk$9���K`�K��4�G��1��i��T�L�+�����'5�Y_�42+D���"D:�� wj^��jA����E��4%�s4�9{4XMs�����Y�AX���XW�L�{V:���>zV�{B<m:<�P��1��0���e�4AM���ӻ�f���ʴ2���̂�(3GY�:oS̈�[�9;�ؐt����H���t�sZya�Ao����� ��R����k���g)T�W�8�RAD��i��w'�z����0>r&V���ww�&���/=�敛*wZ�Jh&n�M�B��
 ��|�"�(���������������2`)J�5�z�k)Z��i�����I�8f�.N	�[�����-�S�#{qb6.���8NY�V���/s�߅��Y,(��;��/X�#Y6�W;-z��sξP� = ���}��ā�8�>7�S�AbxU�ٜ~��n���X�u�Z<Gwe�1�h<'�2���������R�b����&��;�����H�M͢hx�̶ɲ�u.V����7�Q���$�P��'Lf	h4�'�m�K���爸+u�G�b�Ɛ]�w���:tn��(rw���N��r�V��+X��]�*�[�?�|��ę����om�e�:�PG|�Ȳ�����M�K�_�=��Ho��O��%�{�#zN�,�[9���Q��s���Ł�*�Rza@�k9���1yLk�;��i������u,U��I������$�����;�-�H�b�A�2�,;�*�~��\Ѹ��<ō�/���N@�Hɖy !�'Ā/�g��5��A
E��K�T�h�H�I��8��+cD'%����x��Ŭ9s��JL��upKK���*F9�P��~��V��1���Q���d�찌G(�f�k�i�1���Vʀ����KÞИ�o�Z����1��ч����Ѐ7a ����ʋՐO�[�ͳ �]���/��|Nk�o��/�j��t�H,�)a���0�GN��W��s�sV��6-��͡8��O9A6ҋr�W��*�\��G�p&�E�#GL���N�e!�'���1���,C�[��b	6�J��{���S��
�}�.�S<��J w�����eiG4�� ���;cUx�MZ9-��8�u�ܜ�4^��4xy�g�<��/h�5%e��ht�2q�1��5~θc��ե����%��Ċ�e�=���Z=��\v��ߪ}�H�R?�|�l�p� z�``Q/t+���0��WVT�H�h�G�0��e>�����CՅ�{���yg�1���{d�;�_�^E��\Eμ�V�h�x�Ԃ���[�B�D��5:o鯮�QENy'�c���;�W{`�������ƀ���A8�X�
��a�p�{w���B�G�����gz���L� ��H0X�6aƺY�m���D��P�`�B��As��[\�fS6"�s �AuZ����V��?q�O|�]�Pʼ/Q�T<s��]P,N'�es��onq`8%��0�v k���~>���Q_��>��E)��r6����x���K�d�z�#�����}���E�̵�`�
q�k�q@�ZQ�	]$7܏8�`�~�(X`x��˰IAJXA���T��Ю� � ����;��44NvZk��4�^�g�KZ�6��f;�����fUDM��yT��F�|-*�IC����I��+���|~�Dv��6N�ʻ�m$��+M��Q��i�F���u�zS����j�dy���1;z�U�G ��`�Je�
9Գ	o5�A�[J����V�8Ɣ��>��wpT�o�A%Qh�a`�:���UÄ�)���d[w��t����)>Z#@̛E(��G��J[��R��oz(V���c�H��3���G�m���D�f��~��x�TLR���Ƕ�R珅+����xY���tY��
'���,��mҮ��)���z��\��"�x���a�j7���3�����T��s� �]fno��t���^�s�t�N{�\x�R_�i�ץ:~���1����0�K[�JL:>�����\����8��T�,]�?i���/A{��.��,��=�C� ���PB3���:UQ!ɞ��\o���o�W�_�X��(���t��#K��0Kf�x�\�@ů�:RZ��� 4+I2*휜�¿�7��W�O���<���4����`;����Ĥ}!S�~)����Q	a1x��e�|Htc��P6RhB`��`>a�@�0� %\�n~�v�<��t��e�͜'�����׌�->U�WM:Y�oyy�'�#�K���0/R�b�	��v鹚0�|��Qp��%H��:t�`9�~�:TR��B���iW��;8H	yJv���.��h�)���K�0F��i)~Z���r���\���{5V���m�T��VD��^6��n?�r�f�d�E`W*�)���t\uA���^�jֶ�c���RJ
����r�ލ��IaW�cM8�/��R�mMge�K��*1�l(�^�OH_��=���?=�e�K�S��To���U�j����\�J�Z�>���#2o�X�_�]Xη��PR�Fh�5����
(�H�,ѧ���wt��[CN�����TnF_	�ݜ�Vl�oИ���ۥ�r�l���{����!dp��n��=�)o��wˬR��%�U��I���/ir<>Q`��1����Y������S��4�'�*M��)�PE��X �a�=�� Y[�72;F�_)�������ӣW�;���G���~T�An���ԣ/����^�WKR���=��L	����zbe�4d��޶RqX�y���v���	��i�Į	�%a`v�eX�$�,N�7���^�d�	�RVK�8��O�qOT�eҝ�Ne����UPE3�a���١9m��3ٺ��qUR4��iY��M�Aaŧ�)���n��1�d=��m����c�W
҉��`ձQvC�;�i ��4�����-�;u�C��c^l�ؚ=?ETCm��2?`P*R�[��
l6�TI����v�BP�;�xl�9|��yR�C���EK���!WSχ�Z�u�Ȫ&���'�,�K�%�\W�ll4l���Q}�+ ��6����m�7�R?��j����"x�R�Y,"s}A�p��38I{��:�t��I[�}�꼉 ��)��q�sY��t��
I.P̅�
��t��o�(�B���l�Q �Gi$3��
_�<'�[�on.�&� `LB��ͤ*C��bsJx���|�����VVu�y���0�����RVy�w��)f4��Fl#I�۩*��4��,���Q�`�w�C#li��RI�">ȇ/���J���f6�@W7�@����Kn:H����v/;-�(k��T��I�I�m������@�N�����Ss���׬Jyia�n�a��@@���I��(�_N.=|;)�-������W��	�� P�|H��g��5~���vv�66���j�+�J�]X��O��D�E���gq��Qm�^rH�he᭸/�P��
u�"6���&s8>ɔN�~FW��z?Ķ��tK��Z
m'ab��CC�_�C�f^�4�>����'��֦���.�D�Zj,!xt�QD�J7��j��.p�Htc]�v���Yf��n��N�40�����r(�GaLXd~o�]ax��}Q�:Q�`eq�d\χ9M�ǀ�M&�&kyY�֕�n*�����T���P��Mib>;�2�o`�3�>���'�C�u��K�9A�%�oTAx/8�\b�