XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��˺s��Hh��&,�Ɣ([�e%vt�A�|nw�@�>6�E��d�	"��UZ��!��x����u*��S��P�o���]?^��!��y�bv͗�m;,y���e�W�!��4M�á:���Z��ߨ��D�`,�d���{'b�+w�d[�^d�i�F��БO<�����M�5ŵE�u��k���U��	��
��\'�o!�.S�7S�j0FZ�'q�4����w m�U�j��Z �<�1ck'��p��[� ۾;�[��j3��t���g2���wT 5�̻	�If��c1�y���ѻ��D}�oY��$P�m�oʷ�m�yS�;�"�1��̴�����L�O�E��#�COʡ�""�a��Y�=��4f�U�7L�[ÈF!����|��?$�<H���u���*H�
	�sG����˕nF~Ir����ɒ
�f2>O�Vq��h��2�����'Q�48���2�y���ժY��qg�E�gt�K��WNW��FSZ�c:�����9��0O`��=�?�ή�}%���yH3J/6x�3������]��0�z�j&ٖqY�%u�^�w�ې�_x]�ϕ�#�R�\L�ޙ��M�L������b�v��07��p-Q]B���-q���Q�����CD��Ck珊L��.���Hi�o��9W0�ڧ�i;"�y
&L�E�@SP��c���ՠ�0�]pE%�G�9�H�ϡ1�)m�@Eya��]��͢�9 f�Zq���'�B{5�D!�(��XlxVHYEB    1853     810���p��廫��Pj�(
�m���uA-�Nz�S

�qzJ���l�l�y(�����|Luhm�
����`p+����ԁ�//u�V��=I��9T��FA��%Fh�5�����s� uǡ��;y�.���r���|���d��2'q��Vy-�&����	���)��3
΁3_4�E�W'-��Tm��J�yJ��U�\�	R�� �5����+���5>��PL}+D�$NTyk����eU�3[=��4�F=?[��Yh�rK�YB�����uw�I�}��{��R��À�x^J����Wȓ+7�	��ъ�k��s*�7�ʌ�����.]�2�I�0ȩ�!�$S��W�47���$�
�P�Sњ�h�j�<F�V8C-����o�F��'�[I���tZ#�!sܜ�E������E����%�Tȏ�^�G�ۻ�%���]�f}l4���ɾ �#~V�+ee9\���G��$٨Mg����KwsHޢ�^�&�D�
\�gK �,����c�\�*p�]�WuQ�Y�R�J&V���s�:��.�L�����7��L�դ�����G��1����T'ۓuL|��d��44 [C���|̔]#^��f������[��3 �&��˨{AqG(h^����)� ����M�d���O.������1�1t��qV"9�|����AL���:L�ci1�ﾐ�r�f�$��w�iXY�y�4^���%���x��c�-�,�����He��2� ��$�,A��Ē[�gm��Yl~��b=9�R�~d�/1�D��h�H��b�����k�>U�*^�!�ݭ�RqG�E1]i�	X^X�u�w�U���S�;��ؽ�1�	��h�5�mPI
Aîr�f�5ME4jv�� ��{Q��@"������Uh]�#G�3���?I���<�P��ehNL����i��y��K���"��e�i��0���^t�3����%h�|E�t��ě�Վ����wJ�>��Z��BV!`�:� �	)�%`�c��b�b���Y��*�+X,{
��h�! f�2����\�bxG��YiUp�TIFM�<n_Ϣ�Ϝ���@.�jmn���j���^�X)��$����|C�� ��e2��V��J�0=�D�\h�GmdyM��V5/�e�I�՝����b�E��� ��q�ϴv;���a9�w��`W}����e�-�d���+��3E<'��ɕ�@�\t��1�sÀ[����l�Ki=�/.
��^D�Tf�TIX*`���*,�Q<Gv�w�/�,&4' )���(K6��4���HR�U�)l��B�6.�D�R�A�芷o�d�1��w>���t�}usw��B��R���k4�' "�Њf�ݦˣ���Nc~
�-=��I����y\�@{�H�1f=g�5f�Tw�����H�o�sY~G]��k�4��e0���k%�%-���&� �S�2��eXW0�W���%����2��,[g�]������?xnƉ
hW����� �A�<&�m(=�BW@����DÊNh�v�6$/*'�w��&��>״s��NK��|�+�r�����)���u�?v��K9��쌯��O��c��O|�>hfxH?��\���Ț�a
�Ptܪ�6���}����eZ@'�-�����>Z��N����pˇB9Oρp����>>շ�ב�i��D�m�U/�06��֬&�hYR��m}g�%��'�,��I?yG(
���]�yE����tF�od'�T1��9I���z�Wk‍c �C�G!ǵ&�S�팹k�[�E�������V�}�����Wz��a����h������\;ٺ�t0�C��;�����$jk���y��4!�V�e��S��
�a���-��&�/�N�i��{1�Nq�}�žl�I�U�A��yj����0�[b�������ۻ����"j��Q~��U���_s\XX�[{|��@�lI'�a��a���9!�~����I