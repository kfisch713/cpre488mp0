XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���[a�t*���~n�c(OE��fϢ�h�ժ��Ҳ�k<�2�i@]m�<\�*R1�d�}vw��qniJ2��F4kAQ�Ў��������Ua�d;�Ք�����V����,�UjWr�iVI��,4���-g��=�^�=�ۇ��;|!�`+ ����Z�3����9Xl��fau����V���5�`�q(E�@�q4��%�@s�]xp�Vs׃, j=�P�0Y����2V�1���������57���J���So,��]�e��O�iNBq���/�]WD
�NX,�� �^��m��5�'r��r��b�_��*`�sbG�4��9+���f6�l��t��ӊX8�O��E�`˺��d6Gчf�ڀ+��?t�}��-N��r߭�i�<N���ILZ;���	V�`�r(�����r 6-Nc����?[�zib�t�,SL��~]�q��w�	���Y���hf�����6�JX�KB7�[�[�TG>��B
�P���1���do� �1���wD�D��uq'�~x�1��+S\�$Y��e� ˎ���� �0��&��L�8�1!�?규����B��gY|�zK�Ϩ��fN�G�{������FO�݊{�R�xɘh4i1�q�h��D��l��>���z
�oi�b4��U#6��{o5�`������<�����)��)Xǉ+8�>ͤ�]Eۑ4�ds�N��N�;�dzv�+_�H���D���]�"0~����ʎ���_�n�XlxVHYEB    1853     810\a	ގ��,jǴO�Z*�z�g2�P+*�������*U�g��)?�u�ʟ���E4�Xl�e��#���з�V'�u���0Yݟ��������)c����ϒ�Lab�
��G�q�꺷~>��xi�w�����Y����5JF~H�	v�Lħz���gm>�\�i�����D���Z������fo��~uYm����S�(g|<��&D�H�e3[�`�_{_�"=ov��Ig��3h�[�s/�J�nk����t�<#ɟ�B�U^/�ۮ�x�+v�kc�����E�7A��T*�h���L��_��&���u.��<��Q���c��\/������wd�!9�G�)(�Y��.���k�k��4[$y:Nmg)ejd)[�W������	�Z�\��
�U��n[:��^��4.�
FS��-���}�E3��s�	�t��ܪ���7�N����O*��� g���!\��|'���~�{�����>`0l�Z"�)��yWk��&e1D�疌��_�	�E�s�-�Dp^����5�s�)��՘����fv˩`?,�S�`O�	�VU��s?���xBHP��#
#���U$3��$�j�}�U�)�Тh��Q�C#��N���пJ+�e�
���E��+߰"o����^Մ���g���v#E��й��M�3ӗXOd�[�l�,I������J����08���e`���1þ>�qwi%)y�U�ʏ�ӸA���^c<� ?��7�W�i�Q�|����wW�Vl˜��L�F��/��[/��@�f��G�XvX ��z��I�˧l 0O��8!jՙ��S�C�c0�Ռ�9��"��u^[��:��na[q���>@Kk+� �k��S&H������n�
޴�7@��<�L<`�Z�|	�VHiIt�z���KA��{O�<Tk�4��a��]P�Z6������� �HRg�?X�d����I�Бv�;O^���P�ba°�o�u�7�0�T��pm�<���T���hp�4s��M0��e��O���`ARwEeL��R��ֆ�m�Qo����Tlx���B<���^�]������%��Mǃۿ���V�4�q݀%W�F�8����>BM����.�-,��"�v�އ��\�#�8����^�ޔO^{O�+Aݿ��-C��*ʊ2���1AJKh(�Q�-� ���/��|�ujCu3	��PBDGb�my������;g-敻K�Y��ΜO�0�P<�X��6!1�9�`���MQo:���'=���Mv԰�kWR��_l_׿pS���]XF��*��qS���!]>��b��nM;:�e��pr��m&�!��rI�N����9�D��1 ���z�L���]D"�~��LCGZ�KlX/�����lr���w�=mm�z�V�@
�����ՄQwU�8��:�>w�x,�ڙ��2xv����%~n�(K�Ԉ�6KP&,�x�B�D�{��k'64��F]��nw�=�K����xg��wJ��^ݡ{V��s,����nP'Rٜ��W֌:�5Q�	3�:Z����y/4�����1����svx�%� �Ý��yٕ�8D,~���>;�,�n�3��c J��-��jtEMf��'�k�r�K��mҝX�6�4�y7&X�!����'�#�Њ���6:�}�@z���o�F��uAK)�����a|B�HC��j!Y'% =�l�iC��%+��r�ZbeH���Du�^EX���Ѳ������8��hP�?RJ�=%^XRsD{����d�7��O���&y���[��zwZ�M�3o+Yh'��bx���ih^�[��_�[q3��|9���@ͻ&��IY��߼f�5fYZPDb^�cq�.��C��E.ILٕ.����d��xه�ya���	(�*�!G�����]W1�l_���Y+�z��7��п<�␴���d>�Iƃ$QV��*e�b���sP0=�]���"^��s���n5P�<�V��<�g�Za(���,'bLv�7d�!oJ��.J�]�{Ґa�