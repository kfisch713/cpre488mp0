XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���l#TU�����~�$�Ț����s�#I�{;Ѭ��_��H�PT��i����Y� 8����[^Z�7g��Edp>��T��-��ҡ&�G{�HnAg7���o���5���7-0'7:��w�'��y�X�k�
)7�ӊ�aŤ�'�9{s$�!��u1��z�us>|�%��Q��V���&<&)���_I���%B�T���ۚ=�����-3'侨����҄q��a��>�a$���/�`�<�b�+���2G=PhP�S8+�Q(�%��̤�8SL6AmL���+�m�[�;���F��)��,!sL��)�5D�c�%��$d<M�N�Ͼ�>���t m��%Їho
��X�C�X�9<����d���`=���
�L�I�k��#��'��*O�K�s�0��/��3���X������[
g��	����T�o�����e�V�gw2�Y'BgK��R�)�����^2i�&Pb*lo0Z3�q���?u�ș��ZGB`*�y%� �f"5qh����K& 6��a�ϟK���f�E'7!M�dɵ�-�bJ�����s��+ws>�lL�JUy���!<y�F&�_4jxo,>���c�UJ&�, ȻG*�*w2Y=]=���p���S� �f"�.81��/���ȗ��̿��m��BxS�}��6���F�F��V���O9�����f�[mac�ѷ���ϖ�2͛�P��ԩI�q��Xn���/ـ�̒vpEm�SI|�톔�XlxVHYEB    b3c6    25b0{������������J*wޯ�c�� s�� Ҁ��j@e���l�N���R�/�Xc�|ްqsɧ��}���O��01;�h��G��FO��3T�$�D�
{�tS�������e�D/AOW=���b���Rs�[V��9�U�c���@�M�%���7�+�U�GD��0zs*�(X�����ff���5��.j��~����H1����~|l�7*��	�	��=���q����s�gje(�Ӏp�3�\Y��њl��7�	�+uv�:ꛢ8'��`�M��>�����]�����E���Ȓ6sժJL!�23c��xe���b�!3�J�<6��4�jG׫l�`}w������~C�9�t)U��D����S��0yP�)+
��Z.����qٻ�d�LY�ƅ�mSY�I�Ձ���A�І�����h�O�-	#끼 ���5\*F�H�sR�
�)�f�W��1�R�h�#!�d�܄W��
7�Vå�h��/�'r������i�����:��%T ���^p$�`r��+����,>`ް{Ҁ�*,ny󚨳�f�
�r܏>�� ��]E����x�u��`���7�Ӓ����k�jf���R��%����0��W��m�TK�����vpG�x(;�H��7\�K�-��"�)�9��Ç���¾i'Rh{�4��3e�J�ixuy�WČY�3�y�h�f��6V֠�3�_�9E�u4י���4m#s����r~ӺK\8���*�":L�����jR�{�(���9T�Hm9�@	��XU��K'�\��)��E��ʃ��䁻�DC�����ܴ�œﻍv7H%�A�.+��y����sG��w�J���?�z�'�>��������r�c�����k�M�ߴ�P'SH)�=��s]����LK�,A��/���zmS	|e��@�+��Ր��S^kj,��k�:LW��vL��4 �MN=3|�.a��A������_����Å�U����h�B{4��-ߚ؟|�����PԞ0�B�������)�ږ��^Su�X��,T��m��Ҫ=�����6�$&�S�c�W�s�O����ؠa�]�P���n�hQ(��;�wK�v��bY�IW��K}�����>C��
�N�,s"�����(�ڦ9�p�n�I���/�D�����̓����|�Y>�8��Bl�i��~c�H��P���T`��j�`ݶ���~=<S�_���D��_�+�L��B�p��hE@�!¦B%��1�#�^��ZI��lR=�yQ��T�e!�V["����,��j)����1��Up���pc��֠�ФC�����\��l$�s\�m5�F��h�Я1��5�Msx�-�P������T�58�����E8$>R7s_G� ��I��l��g�	Kc̦�B�%U�U��0zw�\�,���}-WCA)�2��u����0�8U5��Z���"�z�*��h���(�e�F��b�B�=ڦb�hҕ�&ؔtMeA����A��r:�M\>Mu$9>Y�P}
��Y���{�P��~�Y�硦H2��������*�&�!���
��>ț��=!� �3�g��*+�\��A�*4N�Ί�� �H(���p	tP��>pU<(�h����Ә*�AZ�R]-@�Em^�8x��w@>3\��[���;3$�[�8�20jf��aj�t��;�s�&�ܵ��oۼ'����x,����P"���ct��ŕ����՝kD����X��9�W��=bP&��6�d��Wy8�%�r�
p̓.�\&|�挪�o�kGS�Q�����n��o����,Ce���<���H�n���.�h��CM�� �Lc�����u��j[�Lh���-����k�>)M�X�Y�������K,o]i����%~y��{ �(>v�(����DJnp2�D�����}S�r��w��3�aB
7ӂ��F�ǂSJG��pitY<�۷Z���II��M�l���F��P7U֋��Սς�n�@�Ur�T����eР����I����bJ���T��H��+���
��m	^y����2C��h��V*`��>/F��5Fk�y�)�Q\1��6*����w��5��i崗�9���Esn%��!�WQU��V�U�$��ڊ�~{dN��*y�Ȁ����Y�U�b���B���2p�z�-�6 A�:@���7��V��B���K~/d���*C"���Z�Wp�P!( �2A���s#{0��V_�/�)�=|X�������Ag�~p��_���������|�����=��>����|�L#�пF�k#~}P�"��VH)�����Y[�Ĉ��3�<v��"D\��V�N��y4���O��¦�t�k������a�B�ߡ����=�Ox�>(��0�t�\�K�����\�~3%'.�j~��hd�!�^h��n����	V	��'�/�t�q��P��,�z<��~L�|�W	Z��/�{�93��Q�枥yL��M�
a��5�0(DVfQ����Gv�ԩ�������	�Vܓ���j1}[�HL���_R��~,/�%����n87�v�ϑ1����mW٨TYr��,�b0?�Bz�x�����$���Zc��MIs����S-IS,�D�����
WI�yJ,$���.��F�q��u�HSUӞ%��C� 8����-T}��7���XW�Rʬ��`7�G�!J�t���&���J��`�<�s��lĵ�5cӑ�-�ͼE���4�]J����gK=���;v/?���V\=RO"�U��ߓv�Q������庹�S�����e�f�S��:���>��d~��ϋ��O�Ӛ���F�1K�T�����k�(Rr:�%�m\�L2�� )�&��3��*�CU����k�����?c�z�;0�P. ��w���6�קHa�c"�[���p����������7Q��WCƮx�"1dR;���\���$Ka�'l=�Sy��0�NT���L,�(���x��Zcr9�>��M�f�Ʉ�+n��쐵u��f�Yc6~i��E�ow�����K��J��i�Lc7�7A���י.��� j��O������(iGr1�U�T��5�(	O~;':�E�s��}�f�x(����˕]Z�E~C���.e�x��j6�����G�n���](|�n��ᔵl���oWV�>"�dG��e�ز��8�]<_��"Q�hf�����0R�}�Ú�t�H<���ғ�(o#��䡼q2�uAxY�	V�ɁD=�7�kh؉kGf����P�_\گi�Z��œ��N�}o���@{ܡ���6,vU��0ɋL����፪B:2��A�~ZBIA8q�ω��#\t�Ĺs�NP����+�.H��NR��Q�)Ӊ	�}^��b��^_g���tho���Fcvyq2A�1@oƬ���w�X�"m7��.���M���U�͹=Ԇ�4U�����մ��t;��	)XN7S�B34d��tG�����-���k������/���ӎd�
-��p zU*^��cM !R^Ù��.���a �� tq��m��_׻V��:L�s�q \��<C��Y�>�e�=�P� @3����#�ZiR˩:��nc/�;��I��5'�3����B�5�T�Y�H�HQ�\�.�s�V՜:O�C�t�F�����3g��c	�@? U�F�_��s��K2u�*W)�,�����m��ص����J����^�G�@��3�]Y�;m{�_��!h�O�)�kt�Y�ﳢ"aE �<΃n��O��h�;��%^�C��� ���������	�z�Z4��a���Ӷ�!��6�[�z��ꤓڅ#���z#�,l x�� ^��"7��w����3�������H.�o��x&��|�d��hg�oe��͵����*����8e3���K�@���ʐ��C��I\ԃ�M���BhLO
�%_�*�k&��������`��� �MZ�A||�����Z����5�JX�0�}*�)j�糠:��f�f���PB�p)Kc��.z{����T�;������ �7�iB$0��O���h,n����C���6F�VP��JR���;(��;�,�j$h���L�]��j��e�w��x�N��Y�w7���p/��>���I"�Q�r��7R��C���E���K�e��y�Ӆ����9$��N=�iT^=כ�c;�j�O��ZP��*���E#z�Z�WNbK1��Fݷ�۝.G�m	�����S��ş�K!x���p����_,�?�c-�Oi�?J�:K3b�!�����9�b���sJ�-:b�N��ݕߖ������5���Г�7�Iǟ��g�;�=ܜH�^s=n���Y]-Jky�&������|}#�R,���P��K��^�VJx<��Ќx��n�*�t?�g~=,��(@?RzA�`!]"�jq��H O������?���4� �yэGg�����gu��CN^�݈����՜���Ώ����WY/�.u�Q�fW�R��耜����[���,���HJ0�C�u����Χ}�@��-�g<���� ��!�\���B������4�a�Q�d^/>��}������ν���[��CȰ�\�ڕ�A���jǷe�U�e��ZΫ1�N��Z0T��F������(^>���f8��Q#৽�X��Dz����+2YW�/J��F�Ȓ�	.��2�(5���p;L�.00�Fi�0O(�+�lI�)�ͪ�W����H�F�#� � �Yw�����"I�f�3pB��E>"湷 �RM5����_�VngF,��!�+g�;��%@���'K�	��� �*!ஹ�@�z`��9�Al�����wHL#���5�ޭ���'Mn�<�����U>e��Ϡ��}ڨ�h��Z��:�K��x���+(�k��:HK�[�����N���Nl�bd��v�\" })�R3�I�%h�u�idu�/APt:d�V�J��`���Xm���,p��2V��\
����ץ+���2��w����$����\\ٶT��G|�.�3��@آ���t1�x�v�;S�G�!��`��H��_9=��f�og��<@�OiY liiZt����*{}��p��F>�l^��nrܠw�� ��'0�Nmr4�@�G��a���Y7��'}�Ӽ�i�Yc*j�\��Yp/�Y���9t�jm�,2z-���V���4����=:!_9#*�SN�Z<�a(2��i���C�飒��;:m��POxt'�U5�1*7�V�B�L����S�M�`ȭj�F���[��Ƿe�h퓆�k����v�(�H�מ��oh�9-+�O%ց��)81h����6�|X�hD��.�$-���z=��LD'�,��Q]���;S?C���e�m��,a]p��r���w����m�t�R�\s�3�غ!�8��u����;��KD�~�~��{�@�j�M�'�����.KuR��~��M��l�/����W�@mS��ؠ(sɜ�c/Wc٩L>��b�OOr�C�w�0��B�\7�w9�y)��r8!�ɱb��ֻ6��E)C���yc]BL�/k�O�p9�k�O������S��	�D�n �	��`��p�P8;-���*�:���R|�ꪸN��J T (|Z]o��х�c�R�e$�[��ʢ�vֵ`!���/N�#�����չ��Hp`	�ȏ�v��^�t�t�����~�L�-��p���3����[��eh}}Y8��ˡ���;��[��q��SS�l]�3n������S�T'G*舴��`p��`Ko_�f�n��Ѯ�R�E��|�{23�c�i�~��'v\�+�Rq��JY��î�wδۑ������[1� �v�} &��وJ%k���"�*Z���O���v��&"�ɳU�>5�ڄ�"ŝp7>>���z�vi��N���N����;-?U���Ê�FK'���m�Y�m	,�|K��e<�c�O(�~�N*�����A;&ո|�Fq�&<rkК��G�X͊����#T��
����{Ng6Ȣ�ȼ 	�C�HGC�������W���=�Y=���S�d�+G y���+�L�J���0���&	����=�M��G���M�6/�	���47�L�,��^����{$v���o����Y������͎�P����Ea(��K��V@�u��,���y��RD��?�k�PXm����܆���Ԋ���.H���%�h�Z�ҝ�a/9��;�WI�j־^�h�{���-�=��cd�a�=gF~�mcJ�fP�"R+<Q�k&ux��r^��_�Z�����G��A� cHp���u�Ň)�rAFp�a�>G�J����fRq)'���_T�?�A���A'I̗�WU:�\���vo1Ҡ�ݼA��6�6#���8�~��Ug�Rp�
_��L���Ȏs�K씭ps+vA�=��)΋y'�����Xu��, L�@�]���E��'���֓�涉�)7{O� �R�z]���<<�%��TP&�uɪ� E\[�V���,S�����IK�:s��>6��юj4@���uǶ8蟌mx�̚Aq9v��Ҽ�#�^}߱�
�VA�)��_�Zo\Y�΢�o�g�.f�<R��*Vr�\��$'ռ0���T��nR#�1�[��-���� ��N A��Ov�;!lV���~� ~u����^N�[�!��"Z%��
�W�@p>�b�1�V��	���X~�yZ5j-^˜�:�\Ul�5w�yl���(u���^�ZK_�B�@DS�@�iE�Cd��2��S�!�աI�����l6�ua�j¿/���ɢ櫀�˧�Dh�p���{Ї�`��l ��-U�-�G}��3��|@W;�������A����$�g�����6b
��
�k��wr=��s�A��͕�g�L*D�����f�oN�.�������PG1����e��d��M��
��9���7����JϬ���@�-1c��b����IQB��&��ˆ��T�����J���kg������Hy��h�r�26��	碲M�dYf�������C�G��˶:��0�V�ʦ���IHH��I������׋N�D�_U,�̣I���;����ȿd[j���ծ��`:��"b̀�T�)'4��E����lKQ���^�����x�����'��ԉ�yh%ْ�`D�fs:���E=�]�S�ue�l�a�H�B|��̺_/�C�߳l�c��t6�N��@4+�p�A���r����M�V`��j�����M�܄[>�<,��M0i}��,����!r�Pvum��Ј��-�G�<�\��r�>vZ�3�0��K��t��#50�z�>g<�9DYǰ�������C*\�?-�R�7K���Qh�����E��I���>�O�Oí�S�j��C],���Z����q.OJԛ�b�?s�Q9���P~i���M�#�:��EK/Wh��5�*>��jp�
��T��
��2��!�2BgHU[���O��U/��ҡ�c���c[��A�xId����LDNg26�76��0ɗ��&"]�K��*�!��	|����qq�g堺�]{K��3�.���Qt���W֫���� sf�y�	w�d��vi�uY�Yk�6�dl�⦴6Vg|�_z��F����Mje{�߾x��&���,{b�M�Y���.�S4�j�����y?���}�Gb�/��M�"�Ll!q/A��:���OQq���WH���`N�<�&%�3�3��V#+g@q㾝@���'g+O恒�/FD�`��l�^c�3�V��D���y�  %�Z�#s}O���xtԃ�OwR|�飝;�J_�y`]/el/�=�����zR���A>jg�;��sw�FO���°�Ê
ભ��=O')'�$�5n�  }Zc�F�`������7��.����Wp��3��γ�+���J��,�̊
��M��f�ؚ�:�HN�HA�GB#"�E�4���g�8�h��d�0*�˓�y��3�ה�º��W-�g�{���#zh�y⇡k1_���+�]_�����%>�3H2�tة1 ����D$LN��n��y���"�A�a*�?�t/�S�7U��|�yݵu1�����n�� �&%L��aUE��{�!|����Y��� ݪ����Ob(�)��������;]ְA�M[��ʬ��oh��1��������a�U���:�.�L �taE��#��R�=�	�x�3�b|��!n�`�* I=e��Z�Jэ���QmT^S�C��:���B�B�Tҁ�v9ۃ��N�jVKО����{��|U�q��P��S�ɳ��:чO*���)Wt�$���V�5^k7#�d����~&`���#@s���0ꓛ��G`���"�9�N��3����y	.����l?���(U�fh�*��d����|�by�⃯0�r8��bQ	+��{�L]�D����.�Y5n
Ȅ�=�+�ȯ�C�ԧa?ͼ�QL؎Sw<Up�q�r�^кp~b\� �F+���l��g�EM�4��!�;LR�E�L�j��_��}6˭)��3��m�qC�DdM.�~��*����������\@-�K�&��$,��z�A����;&�Ol?��)�_l@�ahGo�l�kь�q�d��"g��P��0�9|<�Zy."bG� �o�����<��8(�(���8�/��<�.� ߿�LX���T���)Ԃ�Q��W�g��7�=䦮`�8��¾C'U T�s>��ʰ�P痦��r2�-�D�;�o�LV�Ov���P���.�9�?K!�pw����<>R��4m�9����C���˪Q��1kG>��+Ehu�I�[f���c�~�Mo�NS��n�Z��w�����a�_J�1Ѕ��IO�n�BP������>���G<���B�Ts�M��z��W;9�q��g��Sx�1�@$㹪�g�,�� 6^�Z���]�2-���@��Ǉ��]g�P!*���0�y��Fä	{�����uS˴D\o���jG���\� \���{}�Ѣ�d?�������k���pz�|���$���
[��
]���)W�X݃_k+��&NG5e������C5��'�.���'�L�⢫
���sGq�4l��.�ӻ[��Wj��,BC�BFC�˗˶P�0F�3&��p` ���(�}�F(͒�WQJӘK�+�)�߅ƲR���Xĸ����Og�A���}�0��&����=�&GM�y��P���ͽ*�K���V�+��Ť�ד}��9� �}�R��f`y��k���?z�ꘅ_Chה�"�=�&	�%�V�K�x\��b�θ�u,C-X�U�x��Kd��d�X"�^�1:L*��h�d��}:�!���܋�,H@�!z�?�Kd\8i��:9�o�tZ