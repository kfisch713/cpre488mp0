XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���~*Ȃ�Z���b]e�O��a�˼h��B��B��}�(�D�&C�4��L�Nc֡����txZX��ӷ�,=�v��D?U�ˀH�~�	������p�F�q�d�@'���we?�@�j{�R  s1�<�u1�?���N���ҍ c�"��u��!��/�xi��l?���7,����j/�N��v�s�)�R۝��l��S8����(����w��w��$��X���˲�"�k���S��K��ikj��+�.��Է׍g+��6O�B���0p���nU`�D_��Q8�W���[ ��WRa�ra���s5�r>�w���#�μ7��A�tP����r�Ν���?o����7��d�X�?U���+���*^���\��f}D\G0��hgЕ�~� ��Vq���6C9�w0a���}��,r
��I6�yj�
������D+�����-�^���=����6��/��K3#ƐA.k�7���aտ ���$��*1���с�L�ҍc]�C��
���Rj��:�o���!?������]�:��d���5zD.� �:�A�"����vׅ��ky�㱱��w8��FtB��i��	��V��Q�%{�2� 4�J02&��Nw�aRS��*���#2s�mI����(J�U|\�(�`a�j�E���:o�)7b@@�i
b:� l�ޱ�sc�~�	������$[�n���Q�wQ�����y���$ ���]��Rxa-tt��l+�:����QD��D��8}XlxVHYEB    95d3    18d0=34��h��m�Y�2���y�����c�~�J$ӏ>,��I������P�P�1 C��Q[A���*���WWQ2���i�XJ$8�V@�O�8�U	ɧ㮡*�iWa������g����vv �돐�O����d|�o))���u�P~`�/
�ƫ�s�7��l�m�,?]�>|�?���� 1hEa�X_
�ީ&c1t�c^��AJ��u��B��u�0�(4��c=v	��vR�N㹛� �J�lr���D�ǋ���A˫����1#�?�+�N��
*W.pu��[��N�����r�>a5J[���f|����@�J�~���ï�W <��O��"���%a�D|L�)caa�B���j���^C.��L��r���Y$�Ih��ӃF�h%:�-s�<t=���V��i��;�OM��S0$���1�;z��{Ihm�)Z���>0���=@.J���n��\�5;쮮156-�s�����	F'��f7�q#hd���6N�$�S�"�uu��^�����Dr�*UAn�m!\7���J�/e%FNc%�z��袁��g\���)�c�W�D.af` 8���A��<y�a��`2��M����xL(��s�|�mUʺBJ���萿�Q�_��:�6#��cb܅9A�o¹Q���hq�	Z� $:Đ��pV��ԡ�jB�F$����}��~��Qi(Z�4���P��ZѼ[�n{Ԧ�=�?�Ŋ���w���Ox��0�K?ð�����$�Lk���*+�sb� A�y�Pf��0 ��Ҩ�N�kz
K��Ub�?I��ƭ�v��*�E �U��xN�o�@'�^�us�be�o�ɳ�'?� �2���.h���WM�]a��8�S�2�j�L ��k2/�)ɥ������JVD��)����t���Ǧ0����B&�X���(�6��E0�����EQ���?�B =m�X�}�=�3�y����F�
,J�ө��k;��[= ���]%I ����,���n(�{��<��Aq��������u?��r�;��u������>��������"w��G��7����.1N��B�6��g�e\}Q���S�a�������%,�'� i�T�sw�1ԑkW��@7���a]&WI�O��*�s6R9`���#�2wT�8vB����h뽀G��3`s����\)��)��:t���z1��0D�hl�{OK�n��	;�ۧj�KV�ȿ+�Ab��qC�[�߷� P�q���i3(iZ��r6���Cr����h2iܼ$��h
���dm��j�S�Đ��]�X�l�A����i�/
�*���ƣ���l��v���s`�a?]��O�.����uΊF)��ey.uux�jucH��d�S� ���L�Zgc��ZfH��9��X�&2	���܌�4�p�8�dr��7]/��^��j���"�xN�b�ɽ�[ާ��qL�> X��ݭ�e�%��܋UE�*o��zb0j0~0_��
M��cf�>(�s���;	�b����A�qc)���0 �o'�}��:���_�iOJ�hLu5%d/�]iZ�lI:n��Yh�*���4�����ƙ�i�[,e��I=o�r$Z|�W*
�[#r4i�v����3����JR��Y��7��.��-5#:F���k���}��q�Jy=�����_��y�~ED���s�ǿW��|�mg�OPZn����P���F�;٘yl�_���٩s?]:��|�E���J}h��0�b��q;w
y��à�^t��[��ƶJ�ym��EXQ�p�{ZNa-��'��1v/%&L�N�0��r��Y�O���N|t2�{��3pAI^���#�񘍛Xa��iR��yP��A�oO�̿��/R���K*M�DiB�X���?��ZWT�~M�Q��� �RF�;�Q]W���͍B�%I���em�2�U�	��7/:�@ƹ��u�@%��������/b�/`��l�U�;���$���6��/ĴTiD��{T��Zv�I���N����tӘFn�8!>�_4�m�i�}}u^�iW-��@�a1H�q�$�wi<d��<���wm�n�'��m(~Qė��o�ȣ���+ �t�����O�X���D�k��kmՆ'Wc���.����z|
{L:h+��V �ʢa}��Y�B�2O�D�:1@�o|2��CKAB
h���߄��wGbO���yF�M\� s��E-*oU@_��W�M���==l��%�E������m:G��<P�mG/���\>�)�V;*K�'tv����2_��t�3(�f&|�$#��w�����M�;r��W�E�i���q�P���J�Ϗu�����U倩#t$��A�?Ŵݘ�w�����b�^�o�D�pu�8��0͙���RשV|h����JL���R[��B��(��o�*�C��2��}� ��+`a�w*�/G��3�i6n�Z�k�9(� �^":R�K�R(E�K��Zm��t�s>;	m/B@^tF�7�Z�E_	�s���^��,	u�7YIv~��RV�m��{�m���PS��*~7X|���1��ܽ��(��oc�#���n�=���i������ɲ���l�j�Q���3��r�?6�0;e�����M�׌�J���Ɉ��|W�	ּ{ނ���(���p%�m�`M�ZKM'��v��S����9(���Q�Nk<��'�JA�s{9l���o����]�aof��k�����hA�W͒�a}A8ב(5����A�j�#t��4&n�&Ҁˆ/WRxR��8��m��)8�R�ڨ�d����)���8/�ߑ��2.kJ������Pb�.��C���]P�*�d�&�?!GGVг2�=���2�����~.����&P�i>EKjh�A3�H��ipP�͹�%i�����PG��$�j?��c}�W��������8m7J� g�����i>l�i�M��5����Ǚ]1bv� W�7�ۍf���-�}m��rwS�c��&]�qW�����*��\P�!^�o��,�)�|O;;a�{���w~�!g�O^-9��(�����J�҃5�m�͆���5G=��F~��o������5?��]∛�m��\�����A�p	��W;����uT�@$`~���{��F?\��ނw�e�j)YP􈮬�Lk�\@PgKn1�Ryz�i�*����3}|����/�2`5�DՊ{ �B��޹
�M��p��E�]�:0��M�)�	�w��kS|�H�[h<�8�{*H,���f˅YP�!%�#XYD��IBA?{���U�7ψ��"Rf�@��V������H�E���1\JD}_b��J�k|6��T�*��H)��Z䯡0�n��FL�7�YI���Z�$A'#[w���H��ì����E�F�q��%�U_��?�^j��؞��T�3�T&�i"a���
T��Y�9�_��w���W4$0�m��<i!���Pk,��Ī����O[�U͓4��y#D�9��׹&��e�՞;��l�Gf������W㏯����B�+(.O�\&#L�ޞ�w��p��V]�䍡�r(df-S�h�}���F�N�6G���{]�,e<��×*�G�Ue�$'2���䐿�3\	*��c�b��3��w�MO��>���	���y[�=]�� �i@)`_6�������>S�y���ƔQ0 ��R��Oʎ<e��0t<�)�=�����MG�]z�)��C9�Y��������}<�q=0)�H��I�R�\�.i�6z���E��NoU�z��5���`����=�����}W��Zڵ^}����11�������0�*b�u���֗{�r�'�((�	SLےZ6]�9L������Z����][��E�9nΏ*`'#39U�[`' Y�o����/������~�&�- �3����̄p*�<�
���,?��e_�s��J%�'͟@�>2b1'[Vs�uh�'P���6��3ʙo�}Z��QD <��ٖr�o5�N�C��+���%�M�s)wɥ�Pzq��s �vr��^������r\�]�Q���+~݊�0"�+�o�=����r*�ex�s8�����ci�zS�N܁�N� �Xa��J���u��>�~��Y�۲]J'��r*������J��,�����[Cil,�;��j������\�\�����a�k���H|�A��A��E�5 �˛�7�X�zןc-u�>�}��2dWI(r@���۝r�a)�1��nY���>�P�ވYPN�E0,�9+�9�[Ӏ�� V�,��+s��s��z���X�ұ���ȫ���vu���C��P�H�Y��5��9d���������]n��$�um��zٞV+��y
m�׀��丫�E�\Ǝ�R��Ob�0��o
<d�R2���C[%a"(-]c�&:L�2�|>\�M��*><b��𶞿���b�z5|���d}�!Rq"�I�X���(ܖ�;�DŽb����&�����)Є�+&���vV�y��+c�FǨ̇��L1���l���ShlV(f�P��˗�g���V�(���>i	���硯����b�[��q/��	���>�#i"C. �y���4`�6Ʊ�Y����O�rG��St����X���sς�fF��p�oW����y앀��Ež�l�:���K�}��YD�?���n�v����q�c�^+WWZN㊖�#+P��$�����L�'jN���ַ����5|��^@����}�|�7_^��}[Reu��ZȩP!}:f�f�fFO.�}�Q�eD�[�~���� PY�	�!d=��a�D�R4KaU�+����	ٿ�@;�ٓ�����x��w��co�'Mp�B�����fW�
ו^�A/��Z���N]��9���$F�{����%�'|��j;�I�<5�*m8��;���t���S��iT'��+�ï?--ed�*�Y+V�S�U�
++��3�&|���81�Ӵqj;��gf��y��QÏ���,�
���	�*SV�����������;��h���l�nҷ��i��Zxd� �+!ڗqZ��X��q?d�R�`�j�����40"*�ʖ9R��\h��_?o�r4�N�՛	�yeO�G�M�'!-f�N!.���?�P'0��++�^8�Ŕ7b���_��������br��dI���j�wa�j��I�L2�������\�c��3�0w_M��&S��1M�� ���Ƌ}��rw�#�VӖva����(�#D)Ax@���������VY.�R�c�e%+8<c�_"L�	a��G[v����V���4�b�L�d(K�
�*)\�&�⿰ɺ�Iy�;��u#Xhj毒=t)�Z��Z����b{�Y3{���c��t�P�2^��CݣE͗��\�Q,6���縚[��É��]x�MRi��2�̌cƼ<������U\���R���Y�Qy��ľU��R��~N�Ź��_�Ezn�͟���Y*/��d%kQ�O[�Ya�^#�t�.ɀD[0\n�QX"��=��&q_i�`0��MTH���S�(���m����ڹ����$���x���Ey��p�;���_v3i:?���Y%[L�{��,Z�����6�@�f��۸��)��W\{wf��ⵅ�+�h3m�Վd�s��ǏV��4�����J͇i���[���M��_��� ߕ�)Ji�S�������?���ֽ��' L��Tx�n^?�po�e�Vu�D��@iz���0�U�v��ZɺP��<[�R�^���"q�]��\dSDO��"�U�����V`����o;����Hhу,�����qC�B׽��c���V|M�u���d��i�f|�߁h�xzvN'(��#8 �őD�x���e��h�����r���$L�+_��21�%�}w�ݍ�7���J�ċ�g]��>��B�Poc?�v��&�4���g�R9�@F(�%�Ao�e�TuT�z�	�8|4��[�� +:�Xx�g�f[2��n�au�#�sE���թs�]���������m-Iz��yj�@�k${O.� �[KJo�9ȩ}��A�����Fj�$������3�� �)j��[���d�ݨ������tK0j��t�1��8���T�U�)rt��������-H�)~[��C�6#���7j�k/)�ƣo0�2���_W�