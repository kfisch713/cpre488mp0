XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��q�ј~�P����?#��0*��ٳV4_�G5��h�.�OK�|���`��yyP�Z�����	 �[�8?�{����k��1���}
~��0�,r�1
�����Ox�"f,���܃F�c�4�&��4�"���){|g��R<h���-Z��s�5���Uv�:�� ��2BTįdaq��\1�}�+�<ۛ�,I��^u%hFu����pm��MnK3*+!^W���+�T5�\�X6��*���񟾘Avg�i�-_0G.��0�d�45VhJ49��8!>��]+l�=cԚ���5h��,�^$�:���%�K��6��|/���@c��Wsn�ϗF�ZC�6�he��~���h����3�2d�S�~�����������������,y��;!��M��4(�Q���o6�yrW��JY��}�;g:�]�E|bT$��J|��rVpeT(p���{� �sOC�뭦�]�K�حXo�I�5F�m���I��z��b%�#�&O4_~�=���R.y�w��\eDe'\�m��Z&���C9�x/Y}�����l���'����)Bg�"C�7֟�'b�X�N)��_�	��-Ȟ�V]8�ǀ^������e��ZMr�>�2�Nb��9��?��ez4�}� ��x�Rʹ�;E�c�>����!������Uʳ�����bA�K��#�@2�JV��Ч��)L�.�Mgg�ӕE`�jgB(Gr�u���Ղ�n=I�,��H��XlxVHYEB    6014    1840�aa3��LӘz)(� ��Ys�Y���.r*k]�lCLw[l�B�"}��Њc-L����c�!��=�RV�Hn�B�΋�� �Kg���fʺq�~	6�[�qq�dX�≮��d�#u��nV��JM3�,�V: p��4�j`i)�h���,�-�jی��S��&��ǝC��`i�%�Q�ڑ7�>��m�l��ɓ�n��ݼ�m�;���e|'�8�#��N�w��tO�\v`�r�È~��cԕj�=��~
�q��S�j�d��Z2/n[?���&�t��^�FQq�[F`�]1%ƚj"x���Aj�C���M�}t��mƄ'��]�-2�<A�b���������Q�Y�T�s����q�R[g(�w�'������0~�~&Ӧ53�Cv
a���ș��T��'x��v�v���"������f��������|H�5$��^��\�ah1zI�_�a�o����w��L�J8'���r����:C������j�v�)���$�[i�_�jepD���~�/(�CK�����҂.� �
��uJm��u�b�@^�B�OÁ��F�B�퐶���"n��S�*j��U����B�.����<%��d!���ت�8 ��~��U,)��:�Tbu'ck=�lq�<�x�����-�b*����F#B����lC�@�Q�B�9�a�L�?X��LY�����,B t�CPe��>�<���l����0S�&�KmS^=4.~��䯷!^�z��?%�J�.~�a�)��{�?}�3F�`�UL�e\K��f���E�F����o�dñU��5ldpGcD!1=:��L)S�̳x��Nq#pP�𬆪�:�#P�y�
�'�Y�P�ru�}�7� Xq�gsx��O���~��dQ9���L,��u04�
Fr���yR�U;�j���_�_0��cQ[�I�s�׾뫞AA���J�8��^�vؖA�l��U>n��x�17
	vWu�5/��[E(��P��U����ڻ�Q��P����P��a|��b�juw�9����S�gY�)srUL��ޡ��.Aԕ�<�)b�����
r3����+�s��狀�#�?����6E���̄I��I�w�.�� �v"q�,z���Y�_��8,H�m�5�$sǑC(%|dF�%'り�ĵ�����E�uY%�i�ђgYވmoRd�>P)%�W�@����F�n����[�^���)FJ�'/�e�_
���ы��;�=��C-9;�Jj��=ye ���bѪ�$��ձ�5���g3@��?IB�~{��k��[e&4��>������皲\d���?[a�7�B����{�%��rm�/��Hi�t���z�(Ƕ`���k�9��G��^�_��	�ht�õB3�*ʌc��8�D�W�jl�8��;��{�)7�:O\�/�S��:�55IN@d�6l���L�\�3�M�,��vl��/�;"e?�2�Xؽ�JbN�d�UԻ����2����/���[���w
|�-�SȤ��.7W����׍��J]�QK�#�Wذ�!����50F���Ty}����iHv�L[����g�A�弌��Gj��G<���?���J�J��O�8A����AM��?v|�#�	�I�v.IH5f���&X?�X���PQ�������p�BȪg׫�(��L��׊s�-�� $����(�g������1��i������|��-����r9�P��o��ߠ�l/"��V3�6��-�7!-F2�(��_���t|�W��.T��f�(��Q��R�!4K�.�k>�+c�x�Q�����םZ_pd������Ґ�}&��ބ����E�zB�@��nU�g@��:���dqc���_�i���?id	��^5r���0��Ih�d���j�i�6��֮��H�<N{�1�t�u��?f�����Y���3kē@�X�뤿�̀%9o�����{���{����C��`5���n�s ���՗]�fhJ:�p����b7��dU;�iR�2�l�#4fL�y�$��CkO�,g�|h<��V��������:�Uk�1v�6���s_#F�9��W_��U���s��騀۩ג)�"ۚ�[;|��c��e���q,V�hi`/Tl}��c*���Ǒ�[���ᑤ�C�B�$�fFͨ�-�����h���5k>��<����=���SE�>�����yT����+Q�1�3+Z��?vw���]t��� ާc,N�����@�Wa�$O�,�o��S2��u�ܒcDV���͙��nd�ٮ��i&R=ٟ�ϪsF**�WI^k1���X;|��(�c���J\��lF "��P�(�řKw�(~$2�֢�ǷN82����װi���� ����Ú�^��U�x�?�ˆ 2z���dw���9Л�f�d�x�ᛘн�ub�Ajna ��;�2��/�AU�,�ᅓE�BE�2�v1���O<']����<�ʛt�����l`.2}�i!]{xG�#�)b��03��[�ChR���R�2?x�c|-�>�B�h5������ܗ`�}�0��yY�QV?�.8�}�τ��Ƴִ=�Hg��__��isIyT
|0�t2�>��`7:�7j�w�� ��b!��r����B�����"AQ��@��Y��&m�����Lu�#rr��3���1��4�i��O���@C[&Ng�C�����c�Wc� %�0�Ѕb�^�xp�!�kn���)jE0��8�����������UȒ�@�.�+�PͲ��C�@���a�(��{;F��V�;��l'��HP�;�l�!���B/)�����.�C��:�>ʼ#I�D�h����S��w�^�el��ƻ cc�`N��ÀN�Y����zw���i���h쌅:'Fh�le���ǒ�ɶv�b��F΅ h��m�%K�9Z"�7����s*3~"��������ZY����O�p[���{�ދ��(^�f	Q�Y��|�s��{*�l�\�y���BlzD0�̂�:�M�>�4��Ũ��*�Q�oL�|�1��w�c�x	¾/��7'"�!fSpm�Ȏ�ۥn$,�����_"IBdG��%�1�=����i� xv��M��l���
����Bi�$I�GG�]��u�X�ɧe�5�:����7)�o��n������_U��nd4�����qH��_���ܷA��C���\җ��#-^S,l��%��jV����Q}�@z~f�ɗ'�S���U��be&������(��C	L��g�>ę�ɷ13�8�T�	3h���Q�ԙȭ�UJ�^4�`}rj��m�bTP��=vY�lޝ�n>D*��/�{�(G�f���U�JS�~�Ȕ�|�r�f>_�#lXq�h��7��i����ݵ��w�CΗu���$t�����n�o��W�����ַ2�)�oE���2z�*��&uh�#�.�gӮ���+q��4^�6d˃��:�$���x��)��>�2nHgx�z�ie�ABFԘb����󐡣�Ͱ2q/���[��X?~y�2�G���~
�q�r���S_��RYmҺ���Y��=J�a1�B;QwY7S�-*�����S�A�M���@��7��UAt��gq8=�͝G9J{�Y׶�V��Iz��Ѕ|��baXx;4Pj?�JTْ�Z��-M�kR�=����-�w���&w�wlx2�{�>���搃�'����q\��ry4&7&̣f���D��0y3�h��o��`#�A�l�Y8����%8o���e�O+�G�0:�(�߂���ϻ��^�1V,�	�bKGL��M\���Nl��!��ŉ)�o��p�xÂ��h�8 ��GP�v����⧭T���vT��'���v����� ��Yӻ���?��4+��=N������$�ny6�����Z^5�s������] ���Ş�$9�|�0V�N��n��`Ę|�@BB�d�_�7��ۇ=����v��Vq3p �+�r����W��5?����埲��-��Xe �ߌ��� I�Ͻ��φ�g����I0��<��VMv���re��x��*#9�o�n�r�\=�)r�7����mE�LM}ג�O>+�G`t�, ����� �ad_��'Fs�A�^�2BM�8W�R��ԓMcL�+<w���T�sla���{Q������>m.�gH@�շ�~���4S�p�m��	����˗����P��U�Ȉ,�Y��ל���0���e�-1)���E��A3'�<@-�Y�?ҍ~��U����Y*r�A���Vo��Ӣf����ɘ��w�8!Ț��|�(CB��W�"G�'�eL.�l_�E�mk!0/S��?C�tuk�`��ճ�a��@��Sr�h��Z���Ru�j#�ɵ�9�AQ{�3 2��/I���3N�d�Ĥ�Fn��V��@��7�����e��:\i�6M�o����p)����
�(��P�Y��f?݇�IN�%,�vu�]C]����U�Z1��s�w(F��_$i;Y9�`4����Ж� ��@�Te���n���_����tY�	)�D���_9���.V���1�F@�N�]���Ӵ�_�{Ƽ�a�;�8Z�z;W9OŸNJ�7�mѱ��;���!��a�����`_w�t��E�<־� �R�Q�9@�u�U?��ݿc���w��sR�i=��FO�_����\�ֆ���J�|��������F�H��4v��Q�}��ޓ �P�����֖&HGDT*��֍L�{AR�[�>�h ��*帪���Q8���s,/c��$�~
Tǘ�P����9����=�g�OWM�B����yG���t�co���\hx�Q��Ê��N�7���]3��G�U�:��ԍ�
�L�$�'c��Jέ���Z�Z�t�0 	u��4?���y2�r=�Cl�xg���Ե�62��[z\��;i�T�iX�
���b�}��2V��U(�^B$:�	���2�,]L�ܚ��bx3V�Kt5��V���m<2�C�(��W��\	�BO�r��+�bQ��2�1A�=��΅�����G�h��)5)E�󀤀'@p�f!R��Q����1���i����U옂B�Ɩ9b3���Ζ�Ay���:E�/��D�@PmW��e�L�Gi�u�D7;���`h{�h>�l6��Ʒ��
�yTT:)kn�S9�B!���60��@������j0�1k��c�:�\����Dǿ%F�{��������'�E��$��C�uT�����ޖ�ǋ>�i��Va��(a�`]Zh��]�]��끠��\�A��
��*vR<���ˌ�uzmL�MG��z��Y�\B2�� ���!Yi�T��jL,'��i���������E�`�0��ߍ�$�.������~de�>ć���G���A)2���F�E�����N�GŰ<��x�.�a+,�И�/�j�y�x�����'p�٫DzxT��X��7G{���2N]C)�.����>�h�T�z6�D:@gA%yC{�.��/H��'�}8t��</=�X�"�$��h|6����"�X����'X�e�d�����e^:~-�p;�٘��ς�b�K�ϴ����>C�ۃ��3���:U�yv-����e2gZ�^z���|�A�E{����{�g̸��L]���	qWA���u��y2�^3�I����4x�ɲ��� �넩�M	���@�ØvW����;��i@T��Jo�ƾ�kn�xwe�|�'�C�O`P����%x��6� �|�4U���D�7����Ё�yddR=��b*�P����B8�����ٓ��q��́^�* cj����:˴b^�j���;@E���,n;ґ[J{v�J��g�O�f|K�k^7��
����k�����`Y�tB!U|r7�ƹ������]#��K��>�^��S{�K�*M��Û�e�b��J�ʑkg/���
�saI�'�oˣ���@���Ϩ�L(���s�y�U]0��^p��H�@2I�vv����M����յUHզ����׽�T�