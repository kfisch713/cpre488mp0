XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���̐�7��H�x}���(�Eu`���9 �P'���L[G���b1�Tp$�L]U�[�[�1���_�G{0��wa�7��zY�C3D9-5䂭H�j �~~+�e�@��A���j�t��P�nt���A�<���0�kc�62���r�y�uYbU��:=�1*�7��2���ӑ��wG<���'�l��}z-�,Q��k7�K�"�5�=ہ���o�+S����7��n@�`�l���}�:��5S��8�ŘQ�[t�^���(���5����&��Z2�/����t�"+84��9l91��m������z-6�b��C�,���}�6�%Z�χ�����7��2�Ĝ���-+JX2�O�^{m)7��i4�j@���n��O�H�y����h���R�D�'��<f�ĝCd�	���|(e��#'��ߑ�5�ӥ��?ja��O\��"�	�Wk��n�'���~�G���rl�iQ�odtx���X����ܤ�l�==J�;&���m��P�M�֬
�C���e�E�Rr���?H�j�tL,2:����6�W���$��/���\�� ^��m�&�i:���{G2�8�T�n����n���n���B��
�G�e%s�t]2T47�T�P�Zk"\1C�T�[1� סP3�c|�!7��Y�Pp���|,�[��?��ج��Ƹ�����J����S`�C�愴FC%s��g�!��/1�D�Y?]Y�X��'j���㏳6���J�VXlxVHYEB    fa00    2040
2��L'�ƬH�0�~����
�̏�sL/����?g�|);ǏOs��]r�<4'�����J̀�(0[�����4�T="��.=HpS�A:-F��0|����]����n�+ɝI�<�!;c�OL+\��Wt�9֮z`�YQ��R�I*��ڎ�`QC�޽��r>�Z��悐�O�n��y��ܘ�����u1�䬰��P��q�҆�/3m��.wY���X�1�]AA�������_[2⌴�v��F��iF#��4a���)�^^n�u��(Q<�������myu/Ѝ(�BZ3�X�6�tT �hC@��#�;��+L8�8��ɔ�~	r�[[L��o$ͽҡݔ�&"��v�:},�z?>�v	&�N�����}	�׫}"n���(��b����o�z)�ԓ���r�¼]�d���)���2�<�Hfts3E����:5y�L�V�N3�����Iks�׾�w2DګI��×�C���
�[����!����cM�q������c�I���I)���@����(���b^��>�����(��<Ý8rR0Q�_q�X����Αp�Kr�������ݤ�	:]U��'�0
����4�С�����H��E<������S�C棌}�	�5$tv"NZ8�A5�V٘�����I�bb!��;w�p���B�tܙp6|H�U\"Ӕv^�ZD}�5�g����np+Ȳ�V����c�0_���8lm���!������\�Z��X�I.�Ϯ{|=mc�T|7y7*��Ac�r�Pؾ�J��#�î�Ԛ�'��X&a(�D�&�a�T�<yK�s�$w�)�P�6�	���N�UWL�ƪ]����7��*�+t��t6M�k���џf~.�b_Ex�/�AB�q�>(h$��r��:��aUY����2S�Y#�L����P&�=7gZ����WiS��k�,�uɪQ-b�7ډ�v������9�]��=��)�ۃ�v�^|�O(�
u,����N���1}w�=H�̰&?��?X*J�ʜh.�j�E0u��U�+��Îf��Q�7�g\�/@�����M�|()3��y���x�p����ζ�Ь�*���ϣQ�����R�z&V`����Rj -ģ�����OK]��t�In�N4�lFcx��OhD�^<��'�\D.�bA&�=`w��(�t�ך-�s)ՇC��E!P&�~:^e��\w�I�/.u�6�Ƙ�a�|���{-L�bF�r[���x��u�|���uI�'O�g�7N��l��ʬ�8�5��(C�0Ӏ���t^���-�&���L��_s��-Y�1;�7N�{�S?6��{�	�G�1�qkt���G	N`�!�j�l���O�(��]����Pf5ȴ����4)'{Ə�c�Kc���DgS[����f#�ò���X��pu�K`_������d�^��gB�*\$�Rnߋ$�vRΦr���q���ӄW*�:�"��R�=d���y=;�Ԇr�K6z�K3��ܫ}�Ҷ�9�L�l��Ml��6{��Yn6��:���^Fo:)���H�%c��:�ȼ�M;�ʋ�Ya��/����z�ߘJ���Ң_%�uCl�Hs����km}�X�6�Gz��� ��R�kΊ�[�;���	1�d�����an�?�g�F� 3/v'Zq�D�	w�Iה<��ț{����R��]��Mm��s��'�6K0�_D�NE?���;�����������r��[�)��gQRTm[B��>8����?t�с�>��L��*r�hn;L	H"]�^j΢~s��=�p���׌�e����wOg�Y�,~'�:��T��T���o�������p�z�U���-0����|��SIZr~��5��,�GM�f!k	�jd3gQ,lޘO��8jnr�O����J�?&b���!�o������ݣ��1�DR�鼔w?����$���s���M����W�ƃ�h3w�&��I'p?=���oχ����OU��8lvrnA<�6vl�| ��2<�CV�.ԓ��_��F��x��\��Z�̩Lp�l���h�v:(s��}n�P�]�C}�s�0��h�T8ƙģ-blZ>�$�{�[nz0>Xj{�^�;쩲��H����w���5g�=yT��K´�$�x���5Mݶ$��q5����S@X0S�_~�[��p�'r=�?uK+ߓ�w�cAVX����H�}��#�P�,L��6f6e��01l^*$��g�����&�X��ֽk�Dr��tSGr�k9yxQG�5c]�v�ݹ�A7�O��	80�2&��F8a̤�ɼ�
��[�l�
�N�Ԅ��pg���ԯ���JVJ�Z�%`�|ŏsܓ2���B�)I�F��e?<��ypZ�̳-�e7�<�l�3Ռ�8g��;����m�uU�,C�#��>����/���&/��vs�n爑�<��x�_���,6Z�|MS~?Y�g,\xy��kq�Ax3���p�3��
�XP$Ĺ�7���(;dv�v����HрuG}�s>wbAJ�[������T�lE���ǍH'���
z�����D����O��$��;S$���d���8^�dO/����[#�%���ѷ��x�]ߣ3"N6u��1�)���hEh��� �����`��N�n�h�on��%���N�����&��Z��P�g/ gay4|�%"��4w��T�h笇d:�" �ݣ6Z8���Tn���Xrz��I�J�2��<���Tk��a�"m���_^ӪNx�����=�͕����T�!p��<pH�PLo!�i�]��m9�4��Jtr��:h�#ѫR/�h��U�=�.:�a<$۪�km$�*)��r�����~9۪�m�Pt�в�btE�s��N�I�~��Cr�O�l
h��1(���H5�I-��1c(i�d=��O��B;}�o|�5Z�x�6�i�(DZpy�U�ͫ�v�����^��b�n����5m���C��c�ł�H���dP��1�$u��B(Z2��TK���0�J��%G�Q��X��G�~Fr��"�>��G�ȓk�_S3�U�q����������6��Hj 8)�4��r-~۟��@|w��+#L	^yKB���L��S��x�h�W?��4��9t`Ke�IWJ�He��)!�7�@��,X���	��aj�2*���
Ҏ��DT�N��-T!�����K��Q��#�~Փ"R�l���y��o	f��d�c��b�\�.�s=�{4�o�#��34��I��	(��c|�k�vvO��������C�!4ҩ��!/�2����������.gF��~��q�ދ��f���V�JI?;�]Mc���0P�;��)S^�c*�>�X�
ߦ�"����f�ͻsD<O�f.{�.zwV��y�[mIK��W�ք�IWYЊ(8nkj��E�9�6��0�DA�/�\��Y�� �m�e ;�*V/��ju�q�q����d��Y���?O��=��:����׉�Cw8���7������m��!�GZwe�\�EL5�@Rs-�̣�.m�`m%Ҥ��"HO�N��OǾjw�LQj��,��dlUY�,��CH\�OJ��έۄ��o9���?,�R`�i&_dAL�iCu�_O��=m�[gk#y�	x��uz˷��}1~{��0��ݘ�-��<a�	W�X��k�:SQwAo�}ᯒ��U��<9�|���z����\�77���Zd�˰}C͑0��.іe��A�[R����ζe�ŋ2�6f�*�2Y}?8S案�lenu�^����j�����*;3�&d�F
ă��=��!�J(����n�ro>���=6�<y�8�J����\=��"c���w�(K�}�12��/�5�oX�%btg!�e��i�R:b�e�nf���D
��)Z%��ϋ�9�X�'h���Ə��7�X����
҃��	�23�Ig. _���H9��u�A�B�QtJ.�9t_����w+q!�8�K�м�%>�,�y4�G �>ƌc�Bv�Z�ڹd���9�����R���������}�לe�:�*��4�ڎ��mz^#��lPl��M�ٿ7&�<w|�.키e$����1l���OKJ��`Zq!E�qj�+ř>zF�]/�v��)�,��տV)�XM&8��o�!�槢Z�KP����!!��E�%g�Mux���q[E�����1�NÆ������(ȳGNdY�x׺�w>]�R�ɥy�)f=zLm�-��ǫ۶����P�����G��+���[k�6�%�bK`9q�n��I�l����<��'� �6u���:�a���P+(g���d�h���k�L����?$4oL+��[��q���h�ޱa@ϣA���/��J�^���X��Ţ0K�Y*���ޑA��;���&�	�>��B	��f[l#䥇���1R=�D�pHM�MZ�����L���c���3���X��St$jy�d;�ڪ��c����Y2vx���8���͢�I��%�nD�{;؋_�h��f�W��?v�úq���k���\'(I$S��1��Gu)���J��D�a�`�S�"�����w�ؐ���א��*,wJ��I���y�8���vC�Q�va��98i6:��]�܋���w7
(?�A|��j^&�钌���p���=��K�"&�}� ��$X`;�8.�Z,���VG���������M/�+����<6�6΋�8��+A�|F��џ{2c UU0��trN
l�O�}��P�V_u7tx!�s(ѡ����Ok�˹4�:�����X(�������9��?�j�h;�b���C�$Y��РgH|�?�69v���Huk���ti��=�f���ʗ��/E�O_����@4ߠ�/k{���n=���	h#/-��س]p��^�b�N@�(�a?����p�w_C�o'�>�S���\m�u�/�V0/��$�s%�v�:	�����k2_>�#�;��N������~Z�e̖0�)������L�l�;�ݮh�(�U1��U}K���a#���R�`�4�Zڶ����P`�����2�)j�:����'�m�0/gK�C����%�s~�M�t��M�h�zH�9%up�[5mQ)H]�n����ra��e���������/a�jH�������R&h������:�W�J�#9�h�2��F�,��8�G�7�A^�IP���"q4�Ds���J5kˤk�|��گ��o�5�wq�1��	:�~`|�	x̰��+C��iL8��@�K"k�-�)G��~O��L1e�GEo��_�RDt�!�'vh�M~�vXF�rA^`K�1��3��8�}���{ѩ�J����_�E쑢�|�ۅ2|���ْ2`�\?A��Q(+ ���p�p�|q�i�q8Ta!��$�W�_p[�u��<�� �(�]&�p��{0�Ї��}�(�u�b�' ���,M��t���f���NO��ɇ�.���蛍u��L�!��L'��Y�d2駪����C�`�|r��ԣw����w����I��<�~�qC
J��o��]�H?�)�?�g<p²�*��yh��o��qG���&o���_��'a�B�n�k�}&����WԸrVA*�>�.sʎ4�N�ϡ�gMtի�S:
��:����� p���c�6��~N��re
<^K��.��.@��@��}ڳ#���M��V���X��`�G��H>"e�d��x��?���)}M8�)��������±ti
ÇZ76��� ��(�
����8�8�=͍w��[�ݐ� D:sqa�17��e���� ���L���gbp�q���Ej꫘�~�ֹ��������l�\�kΞ��G�*MnSr����d:S& �[�X�� T+�9c���c�x�.� ��)���V$��}���r��~D�>�W�W��"7�S:����]�qI�\0���N^�O&3�y��{���dn�?pΊ�l��49���>��3\6�g����������c�}mы���*�$�B�.FW��c9~����N����/l"�:�W.T�j 4e��f/4F������V������m7��N������ʋCa:�OݍM)��{���S]TH´C��L�v�ܪx��8p�3�[l�t�)Sp��1���V�H�&�LC��ʌKiV�7S�|!�<^5�_v!��tNY}�KH��h")����. �N�BC�^�i�K�i/��#�3�X�!�6���e:���ްCK8�;/��ǟ�.�s��o��?���rb#�[�90U.9���5y�U	�;�caF�\qU�{�,����z�A�B@�O`�X\�̛^Jx�%��C=��~	�R�xU�v���?y��U�_���/���YI9+<���N��F�!�@D�I���HR��/���,�A���Gx�*;0���
���#)��s�k|`�'��-����No]�&�'���N���r�:���
��K9����W�<�ʤ[U�R\A�l*��jf���`�}5��w|VV��6�S�09�fV�n1 "��!n�X��K��f!����#uӹNj5����Jb�R��]ڊ���]��c��C���5�1D$[9WtH6W��8�E��<���~2�ro�5����9y��W3%%tϏ��`4��\(u�㬩�V"�
���.�����'ĳ��C�|���fqV��]^�O���O�ϟ��<�E�$�pii,�R���ǜ���(a2� t�1�L�_�l'���XU}8m���x7o-��S��{�f�N�Ҥ�wF$C��O�n-�<�P����^���m��ǉ����X|NɃ�?ً��pm;N�b��!NJ� �γ �x�WD�*�&��͕E���j:r��a���0�əS��4��ov�l�)�Y�r�)l*�H*�opX����<�5�LY?LE�~G�S��m���Wd����i�*B���oetF� ����%Nz�܇a#����k�����f���Q�[�
ey]j�v�,8M)�42���tj��
͘��qҞ4/'���|̷��cJ��*̱H�U/�����E�����.`�`w]`�u_ ��w�K�F���ym���x��x��9���2�~R���}���`�*��<���Z�Rkl�@�8�mf��`�˺�xԞ��������ŕ�������O#�6Eh;�bM���}�߁T�8���C9�T*g�*^b&|�U�N�(~U.#J�Ѭ��W��M�6o;��v��X@~ל������>X���v��r�U�� �����b����'`*ͣNX
+�vf%�
���Iu�	aZ�p�
���~I�/����䳢E8�ir�4=�L3�?Č����hX��Qeu�]Sv��5���ɼ���W�o�Qx�i:2ɹ��N���w�64�"Ob�$W�77����7��Szl�n��*��z+h��jf�gVR��dV8�XWT/�eT;+C��`�D����9�i�U�Q<��F 
�H`��� `���MR�i��Y�ZU�=�I^�����4z�C��D�����4�*|��gx6f��0�p�:,��7G��4`�K�I��Q?!#E�w�� 	����x$� ��=ߣ
�Xu>���xB��}��}�B�$	�wDMC��{T�SԻ8F �C���b�0Ԏp�R�E�W&E��\'�Q�ޕ$}��B4 ��J��_4�s�؛���*uQM�?l�d�f#+�£-�O쐸 o䨦MH���G�FW!U'$p��&G���
rɷ�C��1�~r9Dgc���r@W$�S�x;�w�<����*�	�1��=�B*�AN� dL�8�{�Ƅ�h,�����p����6z���J�rVip��&L|�� G�o�v&�(5�Tgі����-�"�
�)H�a��B'G6U�@����/p^�I��\@o��]L����(U΅�6�m���k<zIk��|\s�4+�|2�P�]3*żӪr�)�m�I���P�9 �A�7t���T"��G7���%��wXlxVHYEB    4f62     b50(\~ BIϐ�'����@e�[zC��㣳�)q�Zg���G_��z�Մ��������g��K�G7����G���Q�k)ᬏ�&f��=m�q;�JD1ץށgxP�QD&����Z<?���fX�h��#3_�[����u�r�g���k�	ZD
S� �S��sRRy�L'�)j�
����q�����pv�[t��c*SB ���H+j��薐��0a��K3�S �"�ȱG�s58n��V��iR�x�5�[����ȉ%�ٗ�eq<D4��&[p��^%�zwW_�,���z�kd����\���0�mr
�
mú,r$�$DS����j�L���C�MO]�mH�zE\&'�k��0�@�d�~��zA���`�K���|8�UEVe��`�9��X��D{�~%��)�Pٯ����#U��Ua���F#>eѝ�' �ݘ�2a�������&���{�2��y�|Ͱ8�H9rI��m��k���N��a��H\0*�^Z�3�Ydc�Qgh9�i�XB�K�����(�D]ǟ��*1��A}��1r�	�.���a���F���E���@�8�U�|Yu�p�z0�Q�7���"��wʪ��1�6�2Q,,z��� �U����u^]��˨{����e���P9g�:&���5@��\A��������B*���:Z���<փ� !�L����O}q1�?���8p�� \��V�62��d��֙�:��6�
���W��B>��-����X�݉k,u�������5ܴ��xb��<�E����� y����2X�|����p���#������N��q��P9����ߵ���x�n��kYV��v����8�ow4gx�4��p�hnju�23K�K]A�EZ�X���m���g� ������&vXV<�D���]'�	����]c'7�5�o�!��,B�+��_��kK��"�Q��5A.q��3:�����#a�ke�}����D8�	/PM����hb��{#\jT�'��:����n����'���t�Rl�BK��׊��z���KM�y�����-���8
_�����7l��P��ߟD��.@<J���&����@|W��Q�f�9Wo&��%n̮i��ަ�Q�����;��ˉ�l�2��'�T�*�Oc�b�!���v<���ᅥ�6� "^�GYw��Q�f�VB�C������"��.�M؋"*�CvZ���'��?Q����� ����$B��;%�鿾���wYY#'�)����`�"�!چ���6��[ߚ�2uW])�{k�/�.WWE���^�R���1g��I�Զ�*3���ǿ���Ŵџ�E�7Nv��i�5;֪��sJë��A@n��L�������|�t��v.��>b@��X��c���m"NK0a_�ǦD����~�"NV�g�u	s���E��7��P�p�%6ψ�b��{���g �%�9����J&ć=D��e���{�@�T�BH�Т(�3�7G��s�l��m�.Ҁ1�C�I�	q-��;T�+0�c=�U�<�����<!�D�R���h��Pa�F��y)3G+KJb�`�(�M�Ԙ :�uW�aJ��H%^n�%Sb�=p,Aֺ+�^ti��Ԋ<ȵ�#b�l�;�?0�Di��I��1c��?a�eTZ�}�R����2�_PsZ�ܝ$�H������6�	�@t�Iþ�±��c5o;���"�v^e�/��]>���UKy�}躧���֯�WXC���a�^f��8����/n��茛@�M�)#���z՘Z�O|��}X�q�t�1�V�Cw��J��2�d��K$$��/�7�O�d��,����T�{� 7b����;F�e�$�[������: ~_�Ʋ�o�"��E~�y*0�]�P���uqQT@1Y�����O3$ 5&]Z��u��rc��
V��RY��_�h��κ�궿�H��0*Մ�L?�.�X�2��!6y?0!et:��/�Ӌ�|[p���3�xG�H"+��c\���W�o��OD��9_�"J���w��,�5Һ!q�B�/�ea���/&�y�
D�}���jr�h�MIZ7��i�R�B���r�M�s��)	� ���
Ttwu>�^�����B?��-)�#��sIWL�z�����#	«���N�d�%�}�K���EF�������idgO�}y|b���җ�k�ܦ����1�ǡ �w�M��g6���~�z�_}�(�L�@�H�vlW }yP���!�\$��w���q�H���T�h6�M&>Jk�)����(`�HS�&v�-#�o���v$}g­���I�p���0F:>�D���^���o��s�-�TQx��i����M,�1
��}�pNb�&�;#ִĔ?����Z�ʣ���nU/���&X��Fi��z��Z-�(7��PtH���[���L�%�Lo3�c�ryW-U�o-�����-��Z[ԍP�ה�9�9�T?������.fC�E��Z�Y��u��3g7M�������+<z��g�F#�r��n�v�8�Y-l�&y��'�ĥ�R#x��Wٮ�ܡ·rN��[r�Aa��ݽ9�\�<YO�+N��p��_����cچ9Qm�"f" 1�%A^tWO��0Q�,~s��By�Bk��Q��LY�)�y��7��Y�'}�n7����F]a��v_owه:�Ν@��[��Y��+�j�(�dG����\t�9K��u�Y������s
�꽋ZOF�r@{Y�N(ܭF�@�h6�H��(�#��t6ᨻ��[�
��
it�~K6� �x~��q�\�!��|z�dų��k#�f�
��TT9�{j����	|�#�=��L;�}�?-u�1C