XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��O��S�h���o$��ġv9�o�8{dZ��߾{D~
^����P�����	]�|�������r����m'�s��ý�oU!1�F��D�&�Y#��FɃ?=�Z��,��w�����]I�^��?{s@�[p�Dy��#_��E|�,)8f!#�s�7�-zvب��}/jYݜK�uaD�tʷ 0"��P�{��"�~��f��[�>���r��+1�c}0Pk�MDY%�5���R������X_��gtm�h�U��ˇ� A�A�0nLL��V���6��{��9'��c}%��� `)��[v �����l��M�D � ���\0g�{y��=��#u���ڔ�(�6]�n��/Ü�܃�OMj�MҒ� �xC�j���&P����?<��٦��ǂs[��B��"���� j��)߅ތo��h
�d #����a�ʕ�V�}Z9n,|���Z�����rh�U7�����Z&���ܤ�M�ѨZt�#�3�Ͳy[	�E�C�'��)`�K\�� ÿ%�Q�)K�1�r��D���m��B�z>F��Z�Z�w���w`��M&P�+K���]��_���>�
�,��1���e�o�p�5�q"1�Ν�f��L�P�s����Z�*>�<��T��WF�\�H�p���ܡqȰq
�}���
e��+h�����b%PF���~2`8]&����7P�'�i���,P*��N$>�hs9����Z��y���b�\����܅ʮ�>�XlxVHYEB    6014    1840L��S��9fu#�x��ՏzWJ��D��Vf��m��^����sf+N���E	D57Sg1�:34#�~�<:�i��>��z����T6׈k�[��:���z>)I��8��+��M�I�F<��6i�Z@�{}c[d��1*;V]��u�z��n�"���i��N�"T�=��޵���V��7�\\:Y�ٿ^4UA/�����I��<�C#�E�htvh>�2{[����GÖ���,xۯ���aS�E˹��pp&�<OPW�L *�EB���������A��.�	,�=0t��� (�(��V���$����=�Oz����s������+Y��cf���e��ӧ-f����BEbb ��d�& mq��l�,s��fD�ܐgV�6(#��yiǎ�b�J?4��%�?u�
�5�{"&s��T��3��]��Oڹ�e��%��d7cN�*� �F5k��FVSJ��x���IF�	4f�ov�-A��@��y�1�6�ק�ͪ��Iۚ)��vS�2[��:�.��+��8�|�SJ������|�y@[5F5�뮐1����Yz`w;�{��+e�m��.�Qz��8�NT��`�������.��� �.BB�!$k+\�b����^�t�2Am�6�w;pL�:�DcN��bcxI�1��νZw��`���QQ���^���h^��%q ǟ���(�� $ɺ`	+w��x�"l6(����5������~�P������a@PE%�M�u4�b1|&��pEL3ʃ�2K_�n$v�+�1:n�*�TŌ�d��&����fB����>�X"�U>;��G�.�K��'�������$op�n��¢3 S�U*�M��5���{�[����Z��C�,و}l�t'Ŭ�����i�l�\�|z.���)*VC� c�h�x��HC�7%��k_|�Z,ʿO�6i
�ʈ�79U|����zT���6�������c�g�.BIb��2�@O��A1?;��&_�����.lJ�_�U&!ac�Q����&�Y]����f��g߯�OF�:�8��T��+�
6ZL����|�ahD�mM)�{E<�Mb�ь'�;�ݝ0��c"6d���+����I�{Q�+���V�9u.�n��^	
�d~��6o�OJ�"�#�I�4�|n�{��M>��.��֛�R����ո���
v� ����)z*��n�V,���k+q�mF��p���&�~J�������m&���{���������"�Bo�BԵ�� �L6Ve/���(�1�����T$�JwV�9�C�i=��w��;/�-����w*��.7�N���Zu���I�?����X��e�q�j�M:1�uy'<�
���E{,ǆu��`=�ӥ�ܐ^���&yD�Y r�	��/8A=d������7;o�4Τ�'K!T�-7 �X-����$�:���A�P�Q��MyK3k�ߤ�Ȃ�4�r�'��pm��l$�T�O�X�l6�GK�S��%�]�,0 �O0|8Dc0�i�2��D�H�4�N*$E9ye�&ބ^�/᠏4V�c����>ҭNR�Z��X��<)�M�TN2��P�W�v�.���9d'�5��[J��2e��7H�k�F�/k&�.6�?ͪGl+��6~�A3jժi��h��}�}��? ��zA�M�j�J�����R�&��ÊDp�!G�/�k��5c�KE���,g�'��6+�h��\M7���X�ơ8L�8�r�`h}h߀$/=�(�S����ˤ��%De"��ȚzgWw��ѕ����`����3~<!bm�ÑU!9�"�˖��ZV)J^`����HK//�1#��@�ע�� ֠���A�աx�����/gګ�:n�-�j�R+�2Jm`�&v��D���dG�.!4sK�{iƕ'�P6L�϶��~�������-;�A����&'��S�Qfq\����d��,�9{��j��%�k�GwMjh�Y���
�+PO
�i-�):��l�W�4�,�|8�~)N�M����
'�}yW;*9�������Mz�(��k�� G��~;������&y?�����]U*շ[ȄC������d�:a���
ʷ�i���:{qr�60�{��:�T0X��t(J���j������=�D��¹�rRd��2~#�����#6�0ߴ�ķ�����̍{a�4 ��⠈�Q��=D�g���"J�`�OE�9b���2�ۻ�9:�8��>t\Q�I$>������jǊ����&{�0��z0N̯�NQw������˶��4�+B1q���$ D�tO Mr_D,���?�7�|���N$K/a�����Z5�.����5X�0�%�H^a�\��kwR�~��^����Q���;f��Д%���TIz'������)p]�lV���d�����V5g�>�a��""_=7b:�gi5��HAx��;kE��BU��ܯ9��^�~��k*��&¥�K��7}i>Ċ���X�oi>K������
Tx㍑}�v�D��sT�7}����b�jfi�r��}�y�Я)�Xq����Nwoc��d T�8^G׳(0�$����O�T�뎪/ $$���;#���U?G�����]�M]C��u�RRdp�$2)	V�}��y6�1��K���b�=Ћ?��*����:�t o�ҽ�i����$�ѵ��YFƦ^ $�ŧ��rJ1�٠�g�Q8a/m�j����ײ��Q�YFj��U����a��B �@V;��+[1R�瘥(��O��E>�gk���)�Je�;Z���������ڔ��z��LF����Ӏ��T�'�X���ml�bH���NQ�R.��,[��/B��'�D���.ԌK9&���r����֋y�{��~)0\�.&d�Ky '%[��_���ZD��sLq� �x(���2s�L�P�������wB�����7�E��b����t���r��P:,j��elNѺ��%�c(���l��
`�ۣ �+.#
筂br!�A��?<f2l1�1Ŝf�F�2�;O@��76G��d��KRV7�Z�Qj|u�{̆�@���m��}�W^u0`��"CB́��Yh,9��ݱg�>�q8���GS��V� �������tױ��Ԓ�Q����f�4�c"��ro5�F/�=�$�dF�Z�`R��
�����������ir{�*�5d�!S�ɮ���[�>��"Z ���>��c�	����4r#W��C.�sϏG;ɒ��.��6��Vd��}@�;EHO���	P�8�8p���H�Z�y���t"*��v�2����������_�@���C�p�-.���9�%�E��~q��+|x9�^Է�e���4}\Q��m�~�$yP⾰�� I?i���"�8�lےkU��@hْ�r���ЧK��U�
����a�:�B�n����g(B�0����/Ug�s�EQ�PcjW�*pϤ?�����L�M�g̗J�.���[�0�Ur�{c���QrQg�c�zxb0GN�W�	͢j��R0�A��L�Q���V4����HLp��D�y���;���ag��N��H�VB�E�����ж�BQn UEK+�iy>Z�QB��������xe����m��j5Y�NHE�o��]�BL;���w��
��ҪԊ$]�=�y�D�?.�Q�(�}i���ȡm�"��X�z���]�}[������7S��Ö\mה�TOv:h2��E%'НM���ʼ�VZ���bLi�r}0Gwޗ���r�E�P8�������R������=Z���7��'�W7p��>ƀ��t>��ŉ��0wԏ1 \�?��T"�Q{n�mSb%��ܱ@l�|UF@)��7M���r�w�q�!N$�?�
�����o��.���YJ�@�������
�E��C�iG�x�$w��֧{i� ��t@��䄫7-&��ҳ��:$Lw��g�#<��v(�Pi`/,���E��&U&�'��]����'���DoA6������ؾ�`��B3���B����%ߧ�t_��g�m���uG'Y���ˌƓX��-��L�D��F�.~����TL$E�!E�3���Er���+�\��b�/�.��`3P�o[�C���}C�h
�0.�<,��M��n�FX��B������Zv�F�8(���n�`%y��_6%_��;��.�(*�@������#�F�� ��x��7�ʻ'�s�[C��ߓ��b���4R0��g���GDrV����[,Oj`�i�h���!�|��z�]߹��qn(a�L���C�W�V"`U7@Y9���g��PL�������z�[��T 6X���V����%}���Z�h����wq����U �L�s6�<ܭĿ�"͚���a�V�M��?��)��*Ŗ�7Ɏ�[޺��"�+�%R��}�DY;��Ql���{��4.{����� �!8]CC@�t��F?`��t�ܺ[()�åE�q��dq��?��D�"b3=�}_yw*�%�Ll�#���\4`d_@X��
��2��-�p��W�8�-]K���[="g����Ew�ecp��&D1���d2�Y�X�r�Ό��՚�\�
��P�����	�F> gtyR2�0���T.�4P�����LB��\����}̼U���1�t���A�Õ��!��,�nSy�	�H>b��5ϔ��*&�hָƓ�7�}�q�0F����[՗����{�CW{��¿��:b�j�-����T)�j:�v_�7g�\#Rh���21���l�G�}�ovr4h����@}�~?�n��	�h0z7����i��5���d~pYȏ�EO'��J�
Z0&J����o�6;J�6r,Pm|Py��g�0�F]��I�ys{��8�����1rp�+k:�'9q��K���lc㠡�1y>Ds/aU�t� (�ċ��A
�q�~S8c"��x`NJ�v'�&�����l�?�B��l�I���:��<3�V�)b���S|�]C�QWstxVH������|�uN+�����fx7�=��M?�*�����+a����Rz����Z�W<�GȬ}�Hg1f��(�چ�v�6���B
�}�3'o�Q<�7�R���:��n�y|�e����>/J#�TckC>b�/��S�b��P�*au�ّi��T���Vq���
��|�s��nE�S���|�p1�w`���h'̼5�W���#45�S恿D�W��Ci�r}U�X���+��,���SR*��V*����x
��W�5���%&���-�K��J���q��xN	w�Եz?P�y'bOV�.�|�3��{���u���|�Ы
��x������ &Rfy͑��9a�~H�_��겈�gu,�����O�>�W�i�[���ƘFn\��~㗸W��⧛ڟ��fpb�����pU6w��z���?5i�mQ�w�����g揢�#�	���Q��l4���<%e����ީL�I�y�A��8��߱m�O�>�}��]O풋�W����b�vb�bl`�ty="�,���W���,��w�H����,�z���.��/�bdm�g�8�U��,��8�m���!<� ��nimf��(�,=�چ���J���ӓ�J룅�o{Fp���B���-i���A������[�ķ"��4����㌲�����fX��G��^6�k}9���x�p+���~�9F���S]j<�N	���ֲNsŗ\Â��| `���@:a�}���#}��e��ޙ�+d(�������+/ӒSj?��b��bc�0p��ե�>Q��ygR��o��<���C6���L��Ȣ����oa�0�z�Xu{ݪ�D&�M(��f���͖E��`U�� �엚�Ѱ�? �o*�M�?��5*[�����8P`����J9�x	2���54�����[9~�c�%�����>�?�.S��8���m_mf�/#����r�5���@��ZHO���0q�2c/Z����'��K���L_����{���Z����Ê>��Ğ�#��Pa�@����f�������<�� u�GD��1^�.>���ޢ