XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��!=r:BV�et��XD&"OSۯ���B��� ��Ov�-�\+,m��*��7�.#6vqB׆�J����-�(�(������X. �-�+�"W�!�Ѩ_�߬&�9f},���Y�8Ea���t����O�����{`
>��<G����2�Ӂ�ou�""C1�d�K"�n���g��ʵ]���[	�yǱ�g���̓B��m�Qұ����Y����֊���� g' �029=Yh�9k�V��
��_u;��\��ʖ�Fp��tx�v�գ]�����p5n�٣H#_ԱT�w˛K5�N�"�8<|�hI1�-kU��	2��2͂eg�F{���:>���}�kٻ�������-�~{��K�������%^#�_�*�-M����F�d�m���}x�*!�#�7o��B�BV1�@ ��m��эZ-�%;�mH,�{�i��*p&+U["�Cs�7�uC[?��c�rm,����XD�e_v�V�!�T�;�$�2�+�Ii�w?����h� t0�tfQ�^x���̇��hx�<�Y��NR3����a���ϲ{-��'4M�O�O��*˖SN������3��j�e�9F�ɏy!����_G�@E�XG�ޡ�o �\����R-���S� �ϫ�x��^���3A���~�q�~��d��[��c����cD��X��������5�LDGR�F�r�w�`1p�v6 .0�+^��X����U���!��L�����O(,�R�X6=B�����i�2*�XlxVHYEB    3b09     f80a�ģ��i�[��f�:�L���ʯf��6�Kd��T��*��R��qB�ٽo�_��*��B{�t,�W���!bE�G�B1�V����FѠю������`��E�Y�R~OE�ﮦ�Y����YBtP�.����	T��6����4��^�dR���쯭e�v%�yA:B�ߙ��6~J4!���&r�ӟ���R>����cJZ�u����B�.�ɅsQn,:<�?B����ml���bQ�t�ݷ�pTErهTm�F���զ��G x�f�F~�ۺ����֎�&̼f�~�P������_�7���^���x�J�f��jM>��6���Za���]O�Gg\ vJ�SP?��\�@��+xV�D��R&����s��(^gM�=�f:�z�7t���[!Z�9�f�i��|�ǚn�n|��5s����]��Tߢ�# |?n$*ʆ6�|�HZx����Ź͉�u�>	*�Y�yl-��Z���X<�9�/XA8�����`�������aG�9A�43����c�����W�0e��-���HlC"
E����'�2���X�����Vx���#�B��NXl��eM\5I�@�<����Sp��N��n���� �V���i7��� ㅱ&9$'.eRH��@i��mD.�G��N�c�������]sf}��4�B0-u����j�@"Sv� ����Q²9n����a5���{H$����='�1��)F
��N��/)��{���ĸu(�K�Y�0�)l�xƨ�<ph��� r����5�y��w�$�p�7:Cy�~���C�ˢ_`)���E�}��io��	��o���1��GQ$��ҵ�L����f�\�\����3����o��i�����
;���H����J�~6��aT)��S�z���m�1��SyO?�r�����B�r���ܜ��fٕ���A���\y������m�A����F�m�:��paqE���C+a�2�M�B��J �Y� X<>s�.z��:{�������}�Ji���{��`�����'x����٩{����q�h?��+'Z�&�æ&}.�}� �*3�����3��?�)��:+���`�ʮ��W~TBL�;���BPn�2���O�YY�8��?�PlKf	���I[g� 4[�,'�������?�'��`g����`�p-����ɸy�JM�6����6 ��K�I�b���d���[V;�3���tW:�v�E��͔I̷Z@1* ��վ�ݫ�I-"��+�V�E�y��R#�~bm��]-t�A��.��TM�~a�͆l�!"�v��Ғ`OQ�-��:�����Zݎ����2Ak���[���P�H�_C�U��$�|q��E9�D�7}'yN�� ��El�Tb�/��m�r��#V}/,2ۛ�{4��Բ�`_��$x��ѫ���ʇ���Vr9=��x�M��N.p9�JH�J~���!��M�@���st�/��L�뒰RR�ڠ�� Y�3浗��`<=�,x�Ϛkw��F��d�9��3�([��$Sb+UNՑk)�07|�RLǱ�@K�Յ��t�S=o�GN�� �"챙��׿�Ow��g9� �iĎ$/�u� I���������4�a�����C���xT�>��
u�ecM�CbJa-A��}�b5�Fq�+�'�]��a�<�W˥���i�*���F/�x���	ꆚII�3V.�7�y��`�	�����q�k�
t��K�/<��m`'Fg�XMt�����R5���e�\�>��Ot7ʂ�4x�\����F�w��*������ٵ�N������kG�=G��՜���E9����׵"s~�pw��6CXU�o�I��n���t$c)�D�@��o��dKr�_}� �}p�Q'����Z2�����W�­��f�㏊���kYNIb��LEV��:?G� ����k������g[G���ba��ʮ����G� Z�m���C�b���\������q)<�ZQ�`\i��i2�pE�7sh;�����m��-���8,�?����Ė܎���|"I�Ƨ<�r���/�?%\&f�k�]�t����+J�s��7�̩�İ"�2���]���#�������o�^�3������L+�T���`�k��`HCQ|d��d�8�d1�!��柿�^�p�c嵻g�/-u�D0�|u��XA0��Fs��$w|@ۅ�v�zD{<��?���m��Ü%x�U������y������I�d�����d�k��6�`��g\j�!����]ӷ1#	�p� y4R)m-[F�l �J��^ו��zsq%��;��/�q/���"���E�\)<��l��a��u��z�y�ɽ�J��q=a2��<]3��$Hܸ\X7W~9�6}�"ρe�wi��0�%i�lL��I�r��"��QX�{�ڼY�i�S�l���*��0����y�rZ��笯)��4�i����������j���߸q\(���##�&y�zڜe��5�Ӂ��c��&Ɠ,��m�1I;�o/u�E~��+��h��xxg�}h��1�Ź!'i;Z�Z��	���3=��x���4���:MG��ga�v|���3����4V"�3,ׯ觓D]=T�q1�����۫Y�x�J�R`��sM��y>`�.�
�1ae�$u�nw���#S;����x<�#�Z���Y%���~���d������}y̼����՟�ė\��3᢫2'���R� Tf�S�%]C��	�/�+MTԄWjd[ӭ��%�����+P�Vo�V��U�Ֆ�A�X0Pр�!ȟ����C���9%�r�lD;�����f���S�d�l6��L(R0���9���������'�?^|�%w}�`v6s+�wE�+re*��O��K��@��\��s�
����#2qdqi��.e[Exy�ۊ̼� �\a"G�P���+.1�.�O�HX	����ɺ-��I��6��}|c��,�*>�U���7{��������|�m.n�|G]�粩���I���6�ԓ�~��Χ���z8�]��U4�i!o��[�+��Ǻ��{'h �s}J%.�¸,�\e#C��1ET>EOF���]��g9<�
�6#fEe��\���zin����0�ޫw�aC�i!��8P�-�ټ����.'�S��n�?^��")�^:%I�@�����Lb�����N?t9�a22���T�����P��Tưf|Ե�+�j?�;���#�I�蓡���$?�����&���*3aWcj){�^�2����� a21֞�u���Qxkf�C^]�IG��0 <���}��`}g֌ͣB%RK��p��j�s��*;U��/>��Gʢ��c�,s��̞ �7^�*�<��T��U�og)��q�ܘ�;���P�F��5s�T�.Pq�oylԄ�-c���Ӱ�To/yZT�w~+������ex�N����j���뛹�����Y�^��E��q6x�(�>�	��J;I�<n������Ӻ�a����7B&>?�dd���J��d��,�UN0�IOT�bOM��^������H�}�U�x�Q$� �ީ��U�{�����`�.V��Y�yI@7��C�#3Λ��xV� �Ѥ���4����P���_��Ϯsn��U�+x`F�=��?���$Q+��. U�&��{!�H�qj��:�����`�/��5Us��A�~ݗ������a1%2���?�@���{�a5�iE���o���b���<��-��$��+��l��h�	����I]��4\����Y���(	=q �Z��2o�k�����P�`ٹq������M	1�Ӝ3S�@��Kr�& �8�b��b=��n��䒷��A!�N�x����fT:r笓�� s�