XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D�8�������5�3��f���~F�ȏQ��~w��~�N�f�t�Y!��|j�E�۴h@eʢ�S��Ze���Rc�μ'țl|plp)��VK��q��R�k��B^b^�OO��I���r�j?L�1�����C���a�,��=j����'���H���Tv����o�3_��],���F�3��z��P_�}:���^�rŪ̆C�V�����̝��޴����c(9��-����8\v嚙I0��;[�Ά��6l�U�?�e��@QR<���M�	�sǱ�\�hY2�oź
��$��� Hu,���z*�@[�v{z�R"���.(۾	OzN�A��f1�hq
ϕ�"Ѱ9c;h�>ÈS�2��U�2���� �^.4�� 2n%v^�Lg�Y6G)�B�xU9Mɡ�x�j��(7�o��Ɵ3��L��ё�d]�	�q�ާ#���b/*��a73�R���1k�+O\��σ{fK���3>=�o0��&��1 �@�������vw�*Q�b�?�Ѽ+
f/�tW2ůr���#bq�Xl3tW��z�H�	���;l÷@c8�Ì	�[��˜E�aIL�es���O�>�����9� >`�da�bۘS�g߈I����ޓI��2��'8�M(�	b8�!%�+�]a��X(0��.��0a~�G��x�8f����@���o��@O��y��?�WUӀ��e���,����hha~�Y���T����B�cwu;���Yr$�0�XlxVHYEB    3b09     f80݄[��h|���O�����饣���s&�q4�k�;Ӻ�}�Ɩ_I�f��+"[�c�@����)�A��)Z,8�!*�^��\�\i�{�B�p)E�aO"�k�5#�C��MP?�J���@�ԁ+FO�/�*�-T���C��]�^���:
�N��(7�a=rS0�-����w����Y-��m d�Xu�M�_����0��1��dcd�����,���!�X��_����f5��)�d&��u�]�����:��'XT��k�Uև�� �])m�J�apq ��V-���NP���D������1]IE�|�d�����6�F��}`c�էY���,�<֩�W�9�,l����z�+hHK��9y?�@8��d����5�<��JO���R_=�d�	�jY����t����г�ܰ�#;YV �a �Jxo��_��#�vol��&��ŧU��[C���O
[���p-��2?���"Pt[�����C2�W�]����V1����L�TI��u�D+�>&m��7����
ٞ��S���O@��j<��FAD�D�\Xn,<��*
<a�F#0���`(���$E����q/��}��yܱ�тc�ff�*+�%�o���3z�LFf�l�oX=PV�f�^ce��.L�3u�s�M�0�y�%Q�o+Q��"T2�\��Z
�����)�"��5Nt}$�jU?������3,(�S�j�8���N	V�`I���M��~�pl�����}W�i�e*��_|��L��# Ļ�"��M�3N�#��ts��	Y�\U����Ä��9��^Zp��}�;B��l1g�_��a��8T�@y�d���yF��+�P��z�6�-	�r��zȴ�.G���ץwxܼC%�|�\�X����r8���X�S�\���^��ZJ1~{�^��qc�����&�J/#�6)��u���tʬ9��>f��!���^�a��v����P� 2V��8�Ѝ�j�֔Uf�?�d�N��t��ŵz$�_��RGL�F��V���|pY�z�gv�7`���%X�w��xu�6T�B��^4� �Z想D��p��Φ��0�<��K]�H��4���-k#YsnǓ0�5�UMdW|B�u7��f��v*�閟��:}(�}H�����I�d�S�W(�V�4�Z���Tگ������t��̶�3M�'uC��������`䴣$�1"� �^�Y�q�8fk����`mV=@��lE+SI%L	+��1���l�K�ws/&g4�����^�'\��YoF#89��B&��y�3`Ù��F�:P�u������`�	8i�7�)�a�9YtKa����[�8� �����	�E��o��D���/ ����C��q�_.�6��=K�y��򷞴h��b�қg(W�b�AQ.�悘��;��H����=|��3"�`Fn�)�����|(�NO{.��`�ȶ/��H\M�ay+��J�y���!��>�����ǐn(3�q�,�\ ��}ؑK�-aſP�' C�u.6��W��>Jy�9�k��@U�� {!feK�bGf}�r��\�չ�E��n���|f�1'��E��l]��n�ПT!S�\+��~��VŜ�L���L�a(�d�V�?ށ�4܆)�BOp��\<�!#�.Ǖ�[�3���VDb�`Ż�
G�zK*woiS�'�	� �ed�F6�F,�7�ҵ���J�Y�����Ԃi��ɷ�K�/'ʞ��y�>G��c�sc��0�Z�aؽ1����	@�h�l��5�;�Q����9�ElX�����l�:ի�o���@B4����o�-�=��Y3���(3�ۏ�y��1�����#-��`�01/�Q�L�*�TBI���d�GaEʋ�p������15=�L��o�n3+/��dt�����䞃t�?�i�X+��L�(�z���Q6��u��ض��H�MVؕ6Q|xb��Z+��x�5�?�d���H(�|���P͚ӹff>J�!�.~�o�l̟��Fi-�k!�ig�ϒ� ̀ｚ����Zy}(t�����[�A�dtE�^��&|��Oo�+I��x:�X�֨�#�hL8ڟ�=,Y?��5̍��T��hI7N���f�rN�m9|c�ғГ� :�_���͵w�"b�?-��+HZ��9��>x�,��L�Pc��:�j���(_�AM�K]M����Σº������6���c^��J�l<�=��L�2GgRA��h���o��X�-p���Ԣ�`e�Eiv���Hc^����Rx)��G��X{Nx�K�޻is&Cv�n~�'+���цН��k����-%���(E�?�"Cr��:p��5?(Mv"�A�&�A)M����)�����X��#1���!h<Lꮗ*P1(`�ޞ���b>��e?4m9���("���DmVJ�e�~�1�ӓes�!id�z+k��o&�!hr�P���I;�F�po� ��^֫�	q���89b^�ܟ���os����Y�I+������dX�hΔ��oC!����hMY�N���$�ADp�j��x�.�n]���X2�]�v ����S��&�y]�����A�8��K'�OBg� ���ё'W��gTxf��Włg�S��W��2��ſj�C������_���Nihe�$�E>I=�D�K.q�I�p�͊d)yrX�u�0�7$E�qB�7CĵyK��}���������=���2�)rA�k�~>�Þ�kݳ�p����IBB����E]hN�},�%u�� �^W "!�W��֢�j.��;�if]����m���pr��'���ݫJa�j��}�<77��pҢ�	n�#�
�_>2�n ^4��
�B�^Y�2/�d
���9�E�m� r#v��
jY�5r����v��3pUɵUOƎֱ��%��s�#�"d� ��TIX3|�!��|l0��rIm�έ���`Zv�߹f�Њ�(���s��1�A=���A��Y�Q:�I��'���I�*�4bd�'���r�h�N�l>6�:�6��62F2UW�r�_���N��L���c1d��5l������ɏ*$^#�
S�D�4�G���6�t��'��aw���D'��.K���̰���jK���.�~<�E��w��$��D�Cλs���D�w��r�K��!Oja\b4^>��WQ5�9��o�$�.ߟؐ8^J�$/�Zm���9@���Ǎ�[f!�(2qה	K�]$���}�*�eԀvԫ<��o�^ӌ���`�,�h��O0���іp=E�D�r���!#��9��~�hN�{��Hb:_�{(_U��RC�q�9W2�]���ww\�EĎ.��/J�˝���9�X$}�~���f& G�o*5�ǓaV�s�9T�TH4
�-�����:��?�ݒ�@�^�r�HT0L>RF�s�tM�ɣ��
��@*�qӟ�J�=DR�A���R'�j��v9�χ�r�vSq�"6~�\�̞i�#�Z]������� �dsd�
���3�S���`���
���W��ea��@s�/Bb%��N\w�o�#k�;�n��*�RMe*\��/yй��uT+.�l��&��ԋ`���j�^��,�C�Bs�6m�IÅ`y�kh93\��#q��0�bg��Y?5��I�qH���^��V6f;����fؑFl�Έ4��9����k��/�HWJS[���/$Gy��IM���X2���:F2�ce�h*}�~��P��ߏ)�4��b=H��zF6A��p�����)'U68P�M�-��97%'ѻ����}�;��_z?}��v)����S�[i^x4|w_�w'/o֛,HQ�#���'\��f�5t�ąEM�\	��%9�