XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��]���en8���8a,�
��fӭ�W1���wc�׭���/U$����Q�D��1q����_d6�����m.F�����/�I��+�qx���-�(	@�Nn�L���y���3}�E���]��L�����i��I��sI�^z�Jczon�c�.R�N>ZR�Y�}c�X��t�O�G"�kd���Vo���F�E���e+��a��$�D�ZQ������CՌ �F��B����b�B�Q�f��z0�U�	���c�_�靳|�Վj�<�Q��"�cF�*is�+�;;�4�cN���mC��8C�fiY=�qQ-o�U���J�"�1,>9�;.F�FX�+>d�5B7��٠f��1��q�ԇ�n�q&.�"�lI�,#W���~����*�H�[�.�.r��~�P"L�(ڳS�R�ͩ�׌\��}��M�34��B����
>fQǹ	[�!�mzᶧ�Jw�+�����f�M�:�^)����-"�8O퇗w�[���ZO{�������i�����+�C�)�%��m�H�/�V\WBAg��+A-~"̽Ʉ&!e�b��Q��P�H�3!�6zr:9[�y8����9n����Q�ԹnV�{8V�2A�<��mW�gr��FsX�k25����c����тxRR{�eLQ�Ҵ�`�g�\�gO�����L��P  �{+}͍�x̄���g�9��ưb�b)2�|������c�f��/x�)7B��3��Oސ瀡�O@�#��Y�5;ahj�N��js�Г���XlxVHYEB    3fdc    1160s������C��=&�]ᄖ��NV
�(9�e�t{F'���mA�p���PJh+
�L��xhM�5�]4��r���*[O����9��&��هˏ�����%�*B;VVA$L}�٥��O�s���������ԋ	�y �CV��ͥ���!���ڃwy	4���h��l��sN`�UBms�	*"(x�� �����xz�6���PFNg ��f{���6�H��\��f%���:ȟ��b=jsin��&l-yQ��s)�`����U�L)�=剾㤽����GιӺ���s�m���1Ҽwu�x��MJ�mO�#;j�n|�|6�x�:��&���˅Aqv���P���R�tI���R������*����[�9���`�����>�f�E��~�Qٙ��������mg���"��b��J��������.h����L�j��l�Y'P܇�Ct�[��bZt�,����\r8��?�������g�{�JI�53�ù+�*�ECm�Ʉ�zw��'�G�M~7VϦKL�Y7}�!���(��J��H�W<=ƞ��L1YT���qC�^NL]S��th������38{�%ƌ	�?ⱊ�w���~����l"K�s����U_�
�y6�i�`F�@v��$K:���p�v�J
Fy��)��?�9 ֵ4�%�z�X�@�|�u��'XEZ���@q�'���WʀE4�#a�z�hԭn�B�������j���܌0,̔�F�U?>+G����ER��{�RB�C��O�K#\�0�t&���'��h-��V:X�֮JC���j�f�- un *!.�	�l�^:3p:?��9�yB�1w�+#�S��,;7ʀ�}U����L�G�σ������v ��1'�7��9�ž{r+�Pƃ�wբ]O�Yy�������dO�ȱ�Y�cz�"9~{��k���"!F�� �#�I�ƽP�6�����҈%��*�,�iײ4aY��������^�d�l���bA=�T�\�ls�iM����0��i#�7x�=�"{�г���X��7���=P�S�B]�u�jcM5�W&��J&�@�$Ѫm�!�`^�v����X��`U����d�ʑg�a@����/����RG�M�a� '�],>��É9����!E�jߥ7��g��w�`.Q�W�Ay��o��꟧�>�L��߈a kWeQ��� k���:j�Q�ZZS�L�-$`���vp�I�xX s��[P�b�WZ���PlD M�mߪ���g�1�t�LH�Vˬ:<�U�gn���q���h��TMd�fZ�UѽU�6���:ɱ�A����D�i�tl�lx`W��.u*�6� ��#"&��I��_�y�o�hP��K��3�d^�dmRڇ�],j��`*�/e�/J�ͥ'�ݘ�E!�z��Ż����Ƚ+������\�}����ǡ	�=`Aݔ,������xi�L6�����qks'���Ĳ'� 	��f��j�}�~,� C�>��Z>�*����t�.�XǦIV�=��}̅sPI�I�l�WVD*A�=��F�N�aAʓ1�n�.��*^J������97|�X*uGC�>:.U�ah֙3�QbTI�řJd�������j���?cͰZ�����f��<L��&��E	W��r�Պ+`0��l
����m�.+!d�e��|G;�]u� R�W�P���]�g.�I��T׀ס�Pxe\-7j߬{��!}_b�|���8c4�K�[��  Τ�%� ��{�\vl5i��F^AMZ���O�}�CG6��N8�p�*�� �/��v��6p�-3�Sf�mR)l;��2�mߓ�6��"���_1�p��3Rx���3S��`*/�%0LO�m7�[�!~��)q/T!^\�Q>G>F��]�2r�I� #�ۂ�GCO]q���j7ƣ����#!��:����,�uLm�A���;�ˣ89�����:�:2ꋘ��0S���}�&��'���h=>�{��m�G���%�%���t6	��Mٵ�.���>&ӶZ��&�	�&[I
uKt�6o���)��{��j���R���U�,��֟�ĄvLy�N�]x�f_JJb��U�<2GK��6��a뵶���~�q�?x܌��mgP�mp�T��}��O~�Il)���X{�s��d�$@�rK* Ab������	�ȳ��B���@|�YZ��lZ����]��8���02yr��IV�6�n���˸��������h��I�2!B���VP\t��}�E����m��]e�g���Ql�F~��χ��k�FV�g̠ۻ����LN��b�&�(IbP���@�#����&�����e�����{�qd���������r_ճ`v�,ʹ;�t��Щ�P,��pܽ�݅E?��H���=���Ώ��	��.hvtZHfv?b;�k2}k�|=��`�h�0�#�[��G��DHP�PqRQ�ѐ:A�^K����-�l���2�݋,����W�s^���� ��n���$���)�PA��3%�>�݄@�O�ŝ6P;,��:u�̗��rG7\gtY�U����C��2������~�}��-m�x����c����m~"�v��y� �8�{��֯�*�<��T>��g��'Ju�����!��0�T�=���P��VY���S�A�D�k3�Tߧ<a������m��D�u<�4���}%��5���};7�-I��^л*㎖ؘD��	��̩��ǿNF�Ԍ��bH��{�͌�v����+7_¶�Q#U�i�g�,u),����!G�T��̤�58���^=v���B�b3�ѕɆ�P�H0�C�o�N����}-oK����1����j a�7@�Pa*�E�B����.6�#�?[Ps������V�/�7���B�����f�&FS��X�Z��3l�F�"к[�aF���ׄ��9��A��hf���- ���>?\?�N0��m*�Q�x��I�6�#϶\A�17����ҪN�HwF����D�D�\� �E�th7�J ��s��Q�����#�FY�����.
���\XY27���A]AVm5Y��j����DĻ���.󎭔�+'Pu���^l�lFlC+EK���,[��\Ⱦd�'L���M\H�<s�[ |p2������D-��A��?4w�+
��1R�)�v�*iÂ�_�P'�����\���+��/��,�~�����X�nfÓ�&3:��%��N�,A}f��f ��y�m���*��e���c�M'���0t7/S%��*;�]t!���v��O�g ��ـ��W�*�ZE���XVO}A=�G����]{lзJC��K���|V7���*"A �i�s&����%���\�r�
���.��m>܃�א-2��e�!@	65.����b��X����2ft�qM��8��L��Ik���`?W�@:$��݃p�w�,1G�^�\�Q4:���^�H(���5!�Vy4��v�枕��0�@4f	���H����$�l4��4���&9��j΃��o�P�����9W�����b-�A�l�N��y�F���mu����2�����޴��VX\���Ξ���t�J��֋����)��'�c[�@��c�y�����y۔��,���r���8��g�1��V�Hu��:�k)�OF#]��6�m?eqJ @O}�E��!n�d��mZ~^23"�+,��H�3F7d�6��8>�y�R���J&��@(���sBj֋&���aV��%W`V6ʁD��^��<dk6z��M�a�u@%k�w�����#�:F}Q�d�h����}�����k�����8B���?�F�J�ZQz���l��Խ��F6xu�pV������AJ�4�Jc��w�n��mJO�%� MN�/�%���n�0qU8� sD	g@�j����Q��v��o}׳�C�QY���k��
��
�w4�R�1pݺ�z�!ϧ�G�`=��`�*�Ξh�#��nBXFf�|z'qk�I�����s��Z���ܐ�g�"�ǒb���/��\yl�ZO���MWk���������|�c[\>?}�aX����j�
IN(�ŉ�f�I��������LgD�R�����F��J������o�)�}�6��E��y�����_�b��Db�/ѵ�_x}��@dK��<�r/�Rt���+<���FBϨ�|ǅ�!��X��ܲe��x �N�[YQ'�eKa�Y������)��d����WA�����J�*^ˆBp~����y�MϚ(L�ߐ�˸��!o��sW��)w���h��'� ��
ھ֑��-%�xv���{/߁x�eW=�m['���&xv{Iv�����m{-g��[��}�>��