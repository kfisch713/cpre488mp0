XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���jw�n�JTQ���6W��K7�>�_��K"���A9@�K���t��y�h��R̔6G���Ƿ��za�醕����)�u��/��j 37�uؼ�6.ܸ��<	dϰ�+�|�9?�D�?ﶛi_6����A����?��7L�bg*(�Aߤ���w���l[B	�"��?}�jL������୘9�C@8��d1id��G�O���@�NI=?�dpe���Ŏ���X���Yo��N���XR�H9�Y��WM'���U�}Q�Gj�t���K�C��(�~���N{ߐHlm�=�ur\!�����ˠ�� 44̯�~@7$�V��<Pe:;�oU��7XA�}��|�!/����Tƫۨ�U,a�H��dטP�RCt&9��6�q\�Q���#:�Sb��|w\�$��gѴ*5;g�_�U:�or�k�J���y>e��8"�1m�� ��e���ǧ>�	|��/-�I{��}����o�"O�l��|*�Z�$S�}�H��:�q�t�b��?��<�e�Q�Vp��ό��S�iR�X@n��ї�l�ާ��?��zy3$	qNd�_�e�)K]��/ �1��/j�ښ�Q�毳�V�����%DRAɑP{�z\�!a�Y6`�uj�ض��p��mz�,�:���g��}�V0.�ÖL3�(祏#��^����`��2@�{�����:��P����v:��8.�#�#��	�	�w��]ah��׼��>�H_깫U>���9U��ARC���'����v��XlxVHYEB    95d3    18d0����{��S2GY��x9N�9*(zmY�ګr:��ԓ冱����/�KU6��=Kw��	UF�$(��0�'h���!N[|�S%y�sln����G/�O���L��{s>��?'��ol�i\�x=�Um�q� ���;&������))��U�E!�(���H^��4��!�<0�슣�1Dw�JF+I���@V4|o��`������=:�u �t�D���wh���
�O�����Z���	�}��ǐ-�L���ٲn��.+�h�圪����z�f���I�o��<��DȒ����", �=�覭���и�j�C]xS���]�x���*�*i��U��p��b]9�� �ɦ2���3���j;x���Qǃ#�Z40h
}���Ǭ��2�P��F�)�nHA��o�6��<g���E��Ь��^
�*W*�;ש*u��?�z.�tBu�A�n��}n�_��Dd�Ž�F�釱6E�G�tB-k�I�����u[6�<t�����Fp����6�#I8-_���;
H5��r���(ԍI��mOJsqw"\*�(�`��v�z��`�s�U?;����䌫?}����E��l�=*�ky��� �'z��]�]����3��-���E8QX��r5�ǎH�x�Q0
3J��x�H���L�Ec��m��١hl[���ک[��`��<�j<
��<)�MB�)�DڲjŜ��>d!"hV�j4.=�S�W�IM ����R�j>�$n�ف����K��A�O�@��^+P��ߤ, 3�C54m�� ,�o<�E�!�խ~�`E�HR.;����yo�y��(��%=�p/+꫆_ �!�~�w�pJ��)���0[�y��ž�:Z W�f\���4ښ��������'rZ�N��,�I��t�YK�>�]?vQ,r9��x���&P�aIܫ�<-���cn-��]l-�;u�LX.�EH��6'ѓsi",v��R_�]�����6KS!�'�!_�=��t�f��m�e��z�����+	�\Ȑv"�O�y���o� ��n��Y�:��شC�4�C�ʖ�@��E�2�9G�tz m�_��5�P3��j:RhӢ�9���5����^]�B�����<A`��b2������s&Tg�S,$K�3�\4-f�����F'�S��%k䔖�Y����M䡑pJ���y����SP,%��8�>���B���9�@K{{���T�&�dU����x���!�x�W,g���Ŋ�O/%�X��ʽz���(� 82;$��!�h�B�i/h�B�;ے���� ��X�����'���y?���	$]	�k/�B�R=�$�Xlr����\C��|["�A�{���HA��]_��1RLtƚB��c6�+�n�Czl�f���i2>kϛc ���D���կ�J���7�$�a�P����~�5r�B��Bc��^�(����J�;���c21��ְc�r�+?s�A�5 �#S����E ��� G�j]\�vpIN�r�v��Ҽ�{�C�7�R��C%��e�o&99G�m���1�g����u��k@��������:4l9B�[��!H&�,��x�nL.9�1����\��E�tG'O!������8p|��2f��B�rwf^��������U
��@D��w�6���D�Y�xY��ym8n��3�:�Jn�O�d*��H��+�!�'	���B�e2����qX�d�oDOҐ��s���������O2 %���[�7nB��m�+�V���bD���o�,/�cN���QnT@��wD���Pu]��d��n�U��/��<�h+��`2f���G�Np�2U徣���d��5���43��4	s.�˭�Vu�W8��ߗ3۳� f�-!=��*�~o"�el�&���o��=v�'C9�+ꇌ7�8�!r�LŋS|w0���g pL߀l�~h�ɵ8�(uO�&_��K�m����e�T2��3o�d�~��18]�������W��}A�y')@2�vA���	�X�\7G��h,t�/��h��_[w���`+Z�T���%��f���]���kC Sª�)�'��ҪD�Dl�N��@���r>�O�{Z��@��z��Z�U\���@�� �3�K���4z��t�L>r;�����d(��P�P�T����9�%��5�-P�Beq<RG���7QZ�A���CK7���BC�%&>X=ΚS�u�������1���@O>{|L�x̳��;��h��#:\�|�#��0kK=7u(��!k�j�%	�.S�v�sz<�A���ث/RM�__�`֩�Ԟ��vu�uj��o��|��=�C�@��U:��ęH4	��t�J�>B��p7��U�L�n-�d"���+=oTlG���^(����D�=;�������F���@�=5N�ِ���¶2�ܰ��e��ܵwY*� ��</�� "d7���)<K��t߮W�HW�7b0JNf�ĥ<f|y�%�q�����D��5� =!�<���8kc���p�/5M�:�3??F���̎�n+�B�������W�ps��Q��3�XѸ�zy��O:(�`�Į�	zW��
���[i7���u|�LP�h��(��%9,�
�e e�F��� rC/�s�K�ra�c�~�Rc@���#+��ě-��C,?g�,�GH)j�IW8�*�����qum���U'3�3�J6|��ً���)�R����gL�똍�[�IL���X�n��S��c���+f�dF?g86<-f��7Iqj�j�8|����&��y�����,�꠽�����@�ԃ���Q��cWj(���e������^����t«����p d=F8�t��d`#������r�E���y!�Ħ�ɩM�y{�M��'7"�����X*Pf�2��Q �}'f~.vs/-�$���]6�a#i7��;':��|ٌ�]����	\�M`��Q`�Q"c-ڡ���ܶg���*�EM
���<��y���~M/"ƒf�*4w�x�����K���Y���CPG����������Q��)1��E~ ��
��Üu�����̈J�'M�W��dk�B*<骝f6�c�}��4��9���꽰	E�h���$G���A}�N㟰�mm�����~;��QmQ���ω�����z:�h��u^�w`;�Hx3q��N�f�O$�j�H.��>��t��8�w�ե	�1�h����M�f�'*h�Tr[�5z���WG*��Ց�w�g��j��N�vǃ�ٝ.���j0_k}��X7`z8��eB-�O�kd�#���
nS��,�
ǝ�
�<2 �~���d��#��:A��.�Y���(z��P<�� N=U�?�CRc|�.S��K��d��x�A�|� �ry���f�i@�i�k9<����-7�GQ��Ae�+%��Y>��s��Q�;��Q��(���(��Ѱ�W�ޫ���r)�8{�N�;�DE�i�\���n�N�fÇ<�-q䣍BO��(�'����t����Uc���b��F7% �K<�v3Y^�W�.����$���

��j���^�0�_M{A��$��JH ��]0\��T� ,���` i�U��oe�8�����Wiഹ���Y�#�]�A/�67n��#�)��Ǳ&��U�\&��u�/�Ϻ��@�Dw�:K(�pc����tLv*G_Ri��!��������W�Ͻ˚���,iq�1A��΃��JՙF1�*���bZa��+��k@�
ۮ�e���s<��KKu�Fk�UI+�A�oWr��^sA�K��+Y �ꆋ�[[< �z�M
�Гgv8g<X��2eK�\'��e~�?�Z�ƳY��f�MQ� ���H�62���@q�&O-��t��z�у��k��Z=3�<��ݰ>k���;	p�xc^>��~�i#�P&�#b���E�P�ծD
/'؁�ʭ
�m��YI�+�O�'[����a����\����&t�M�*�\��qzy #�k��ǅ�4X݄�lF��Z�fL9ac�͊��'� �Q��&�X��LJ�VV9v��;����v�N(2P�["�L���!��tE��A����@�����/�ȷ���ע��;m�9@Dn� �,�����ze��-�X�j�Q�� �ԘՉ�6���`�VMT��`�9�\ q����/���^��Ֆ�LڴAM��'��|$�!�@� (tW���A�ou]Ƽ�4��[���^!��P]5ξ��d:��.\�GR�R����N6�q�n�J�w�	��].����Ca�$�អ�-Q�!A��~)L%�H*�P����<�?��Z������*������LS]JI�h�w��g�yҍ�i���Ry�	�g��r��bJ�:�2���'��~�4�6:�W �҃y��;��Z�mUQGخ'�,I6�2� ��3�� �D�m��Y�B�uhO�*ɢ��p��j̇-=J�Q�"��f�W�)1�T���~�����7�gKjF�Hl��%ϺИEOEx�c�@閟�R�ll����?"�����q-�&�����w���	����d��y�|l�Ԋ7�I�\�oѕ{#�9V1ٿ�V�$N�ܺ��ѨG�>@�#eVke��U�X
�_9i�]�Bޢ���&H-�}��A�M��<F��i�fmH"O��*q[r�Bxֺd۶-f���hБW���#���,����`��O��%/����q*=������$/��d�����6���N�s��k w*l��0<�H9�𻌦s�zPX�����c���	�/_�N��(7(6�dp5�g�y��1T�5��wت�M����s��Q��$�N��!�c��d��G:0��,�F,��ۆ˝*0��~bڭ(Q�]���g ݒ�pTn�;��1v��G���{z��P��N�]�P�u�p3��a�;`��Y����j$Z�.R���w�(ْ' �&ֈ���ƈ���5g��W(����A7礏�.,�|�s	�H�Vj�!ęE�	e�W��".�ǔ=T�lY�O��Մ	�`�y(�%Lu4�W�"C�J���I��aOUƎR�����Oy�5ѽ_xhR��ΙW������G��_]�?\�17Y�0N$'?���{�h� =�(����}#��?��3�~�C]�J�	|h�H�%s��(x�LE�M��L�M"]�v�f��h�4UK�ɩ&I�ֳ�ig�7yWj��<�쾹] e�s^K5��_�C�Y0Q��7oJW��;������/�Mi�Jt�Xn�î�=A���bT6<5-�n�8���t,A��$�2Ӑ�\&���>����и�<^����
���7ac�+:��K��n�I��"(n��A�2y��Dx��}˥D�=	���tW�%�Nx<���T0:�hs{�ܩ!��W���X%�wBط,?u+�f���o��:6p����ZH,��ϻż���z-/�TQWq��l��e��F��IX�~�o��I�<�8���|R	���(g4��r�d�����y���B�5s'�X�N"t�\�JT�91�W�S<��U=� 3�xyz��J�L6E�2)2�.��˯ދ/�,�����s�Tl���_~@+ijS÷H��j-DHQ��s����'�1C�ţ,��Z�D7EZ5`}f��.׈�$PW����O���M!v`e�甗h�-�@�˙H���6�Q73�r�$M�H_�oe���I�y���+���Rzي?�'��ݞ@oܹ�{`>��y};t
jX�۪b�=�P����o�Gσ@�h��,׉ɡ���X��β�-ZK���{�����kF�Ы��s},AWu0㻺+�!��ěx}|	k��u�����û�3JIH!9V��.�O�cr}�Q�*���F�A�F�� �����Ӫu�@[��9�,1��8O@#G�7����U�y`ڙ���m���[�B�y��:�r$�-���G��m��<���Gh_`f�}$A@���i��g�RϾ_��Df$~37�y�!��w�ы'��՟6p���|ȿk��*'�8Z��L��]J7Y�T�>�+QvS�V�5��%�������4	5N���Kx#>(���B�ָ�@�}��J8�Ǧ��a
�+�O}��^�����)��N��gdcH����,#<0��t�L0g�t��� �K�NZA �Ĩ��.��Z����0&�L��C�F����