XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Q��c���(�:q&��Ϗy7��(.<���%�1��h�u\F��s	�ȶ}��ؼ��2�f�����-���u��JEބΌ˗���6�䳪�vSr,�V��|���Q�99s�*�~�q�lR�y��)4Ǎ�jx;'~��YWjj����a	��X��QL�����*�xleD`�.�����Nl-��<y+�R:x
`硛a�bE��_�'�c��G�x�	���oQ^3� )�!�^o�dn0�n�|��〦N�Tu`g���V~�I��~<T�WDk�	���gT��[��1����� �
h��<%�߁lU(H:2�������(���S�xW��ː�#c(ԋ~%��x�]U�G"�Yzs�X���Х��^|���m���E����m�ԃ+����y�4uǊ�'5.ՏU����A���3١�	�vv9h�%&;й�^]��,�x�EM��s=`��B;�Gfw�S^`�^�9��L�5h�a+�k(Ԣc��#�
7�͌�"J].��	��x�Fg��䍱���"-����ߡ?%�+�ѱ&�^�5�߂]��!����e��&����-e���r/�8׿�;g�~+�w?�3�8��k���h����1�]��=�� �=A�J<�T�&��.�g���.���휄��~t��Q'y5���Eԓ��G$0�b�Ţn����Ǉ_WԈ]�dʖT�%�_�8tS� Pvoh��Ĩܲ,�(�V,�X��DL� ϴ��5���c����8�̡�D�XlxVHYEB    fa00    2040 �S-�PA� ��I�3Ѭ��>/C��4��=�;�>t\�+�V�G��0�R(�Zє׮�ʗI��cS������K���_h�Wt�|�D�P'
�J\s(�T�F�����)��%qFĝ�TD��C㺥)V:ą�A�"�n�w�� p��2�	�{�$*F2�(q�<O��N\�vD<)X�kN��sݍ(����m�ij$�Ϻ���^�I���	&�1��b�6AF�h¶�W�:*j�PZ��*06�`�	)o�m�EM�1},EHʲ�#���O���x�n|�Z��վM_(�:%��S�0ćI�D�S���3��Z]�}��7{�)垏 �B�?��������L�D3�Ԛwn�џ�-����� N���>���`o��%Q�qnG,���q��{d�$AF����v��ii�/+�������]��;Y�/\V;b��r(���-�T>�`mFk=@�|l̩Н�0%O�j9~�+qg����&��Y~_z,k��?萃��1ko�/����%�(L��	�!��"H#4����e���k�Hf�s�
�3v( ��b�m���%�*�.G�y/4/͡?St.ShIɕ�PB����I~1&8�gE\�&dFr�E[>N�&�A�b�u�u��� Y���e����k�>&f���@���n�0ڏ�Z�o�WMcb�!
!t��a~�ż�@��?��&�*͹ўp�����"�a��X�Z��{���Q�r^'��X�۱Y>ˡ���gmĪ�F�+����ՖY`�!���aT������tD#��=:�qt�=��ù�w��uNd�_0ڋ%����L����(-[�ŉ/nX9GLΡ
���m7�7�����B}f4��{���v��'&X
�L�F�3d Ã�D,"���4�����BR@���G�g2a׍ی����DH�ʊ�h��?d���q����io���`W:Hu�o��h��m``yO@��et��Ŭ}7��ў>�&�:t�B�jo�\������3GS�+��\\-P�ܭ���󡋱H�eˌ�e�|�-��ڌ2ikP%X̸�t�w<�yi�Au�����d��`�����I�%7�1�qun�a��f�y�2��Td]"�z�b��5O�~m�	��_�7ߜ��'`�w�4�~Y���C��K�_��>PԸYĠ���L9��(`z)t���"����0�����[>ڠR�3���߫��BM�!���-U�� 0p����'WyG����o0���� V�,iF�������@f���T��0�,�y�6G��y�Z
��?<��G�f�^L�����@� �y�qq����K�� �ҿ�pe��j��y�x�^���7jWLW3-�1��j�ib�I�W���e���_R���	#�0GS��K�%'����S��=���fmO$��˒��.3X�LC�r�5,��[�E��Ky��ר���J@��E5η^P9���(&����5�c=���N��1����=�w��1D���A	GO�"}D@fo���0u��w�E����QD�I'y��-CͧHIRo��x�$9<��I���@�YFz�.s0&�܅��l��U���8�B�R+��W�Q�$r�d�`>�w�~��٢��j}7iAi����S�S��s�|����O��&�"�oa��H�/9�yV_Q�Q��F���&f��eB?�N����w��v}���SG�
��س��x�|[	����Ip�nӷq�UP�� �,��R�uDa��R2�f��#򪅄�m�6\�CJiͯ}���z��ω+��}��:�g�<��bHc�d7�	��Á���3�2��W�mj���mx�N�:\^`%�����a�?q��`d^�4��Y�Z���:�x���$e�k�'Ye����M��>�+XTg����RHc牱����RD�����ַ�%�1���.���������|P!00Bve���B�� �u'꾳������N�I���j� ��GZf���Ą�K�)R�����k�쳄�;F�W�j���A�<��j �a8�h�=�ny�XdW��h�R�Z�ݒ�i����݃�o��;L٤r��сfTX~DT�6��0�B<.B��4�O�9g�j"��/�:t�1��X�،����h�[��i�1:M:R���F+�5��G �K�>`SX����r�n!���	eK�?�{a�Y)Fmwh|ʋt���\ܼ
%��a��f�����`2j�A�\�Ћ1�	(�$&����]y�����Ff�qs�%'��גyy�:)|�=�nd�J�U��;�M��ݠM3�62s�R#�����y�r��\;o;�H:R�2@M���)��	R��V��K��a��@�pLd�N�*
ɯC	��)s���W*��u��2,�W}�׀����S�����2���F�Ӯ8�T�ײ��i�ŵ2C���`����O���_O�MP�_�"ΐ�N�q��u��s��!��>S�J%�Hc/9��	_��������s΀}������>S�W�-m�O�zG�����^%�	ɴO��i[Bg+��=�ߞ������kÐ�DϷ�r{����M�����L(��j��(_��w�}ż�����(RL#R��q���.$.�b�q��tB�8�缿��ׇ�Ww�I�d���iZ����)#��/���2��46����L�߫	�u:� ��8Q>���w�$���a&�+����^F�V�$���`�Ë�(*�Ѣ�!,�*��B���x#�& �<�D��b��:;���E�����"��RZ �QJ�wOx���8oC��q��[�/#�>��CΛ!��Y�!!1�H^W��wPrQ-��̈́��*C��k��������¾^-,�R��Y��ÃN��㡉ш��X��gG)G^��8Y��^��T��L��Ϸօ�����#�gb5R�{��0h �Xj�E%�N�q2O��K[	� v�
�ԧN.R�kׁ^��"���#�ni�<�JY,'��5L��D1R i6SA��1WU�M�Õ�)�(^O���2�+&�+T���E9Q�_�w�&$5N��b�l���a�q��魤����P��D������"ܜ��{v~�-s�vxinZ^g[�B���hl��^�&K�et��0m3��( �iO���ўJ�l{1��Q���߫����ȁ(����fO�&� ��xB�G�_|�W���ڢ��/m��L* όB)J���-�aku�x�n�i܁[��F�f1�3��#/��^A���{o�gL5Lu���uOD�<����/��4���S���a*!�5Wg\���'��<UjQ�u�� SP�R�m�S�^�W���-��,�k{�s�/;c��@ _�%�H���� ?q�#D�sc����9�`��[��7G�wN��֢,V[���5*�!߁Y�\ i�Ɏ(�/�0�{f�dB�>OL���w�az�
Cb �����W!��$�P[���[��K�e~�����g�������t���#�Q"�7G{�h���ZV�Pڠ��������7|��I'-��O�q,�dQI�?s�K���l�L5���Ezq��wRs��Ʃ�іG\�o�Q�:��2@�?`:�r�-�!�z��� K�����l��������o=*�@*���犯W��E�!E!G�g/��Fj�~����%�<oB����}��{)�����F�J�-����'�h` ����zN����UE�ۏ���!�W�cˤ<���J&|�%x�*��CWU��١�>Rv��Hf�:?���q
aD>�
I�� �s�4{֦0}���>[f�V�S_�HO������n�Pa�W�N�9�T��ԭXb��k�e�	��Bk�Yς8�*v�vJ��1J w�̿;èI8���8S��9c�75Vd@T�k��3���_t"�h7CƯ��T�v��Y㏏uS=%,@�Te_H����M�B��^x"��M{e�w�#��/�B/��{�Z0Z�ʡP�|���ƪ08����+B���N��<�<�Fk �UV����IT��,�ߨ{
�B�|U*�Em��*X�u�F�_~/�����7�VDLD�yBv�t���Z�\��L�k]���@Ԣ�ι6$�&%�K5jж��u�rl)|�k�P�)��#���$M��M���(zzl�-.d�@�M�}а\�-����ݸ��0� ���-�һ�-�8~64�r��������*83��S?͂ǑY<
c�
 ��pы<X�=�TZ#*����,H�*�'0�
"Q�hy�x4��>�F��
=Id4�i��݅��Q0]�?(�&ᖄS�.��U�L7vt1���%']�FA�lG��7���Ԣ�����QN�JzٜB��X,����]_J���2; �TO/�CЬ�=z��y��l�~Oy�'�28p�)!�V�9)B�K�[  �˖�][E���涎.y���-Xw�5�i!!����ͩg�P�S�Xl�8���^On�������E��p��sN����h
�:��[��%MI=�tܖ�5���Ԛ(����1�e�-��D_]}����k�-_��(���q�럢���O�ʳ/֥PZ��S�X�f�|?�;�ӱd�?�\o�R�(#W�\Ef����q�Q�t�=	����[Ӏ�]��	{�oO���b�e.�gX!�t�GW.Q��s6f���gJ��bd�y�<%0|�%�}Q�m�ts>E,�<>�9Y�j$����2PP��!�S�t
�iO�u\�:����dh�Q���
WW�xQS�lm��췭9����ϰB�)3��a���te�n#��d��#��P;%g�-�Znhlq���.���W��p����'�u�'��d�����g�M��U{� �e�rm{��?k�,�"׸znrwFQ�[���Y�'+oxZ,Ca� �O�{��U�:i+�ɷWz��c�a��L�E�1�
:��3:�Ԏc��v/K�A�"�'���p�)�۷َ�V�w��v�w�����|�	%�kA!@�ܾ��<�pc�|���Ĕ���v� �F���w�9�>$CH�՛��=�6���u���B�1�Яw%I���K7�dx��2��0؀z~��ǖH7/�a1s�ͮKK�5L&
� � k�p��p�i��`�!גʈ����=]}�B���Y����s�ܽ��Nh�Ƈ�K+�PF��H9k݌A|��Ē�4��K��.4�R| vE��\��ԉ��p��-,!���ǳ���2��v�:�CǇ�~*�l� k,���m�78l���2�?�}��Lm�j�*��c���oU���F�澏��)�i7����Ω���O�]�CH�ͱ��}�m"���<���8Í���Df�p�V=�vvFq���]�̟�tL�u8#��H#�_�v�?)Z5�gG�x�$L�����-���+������M�ή}T.�A8�g�O�9�G�&�:ɤ̫�@��L���!�Gɍ{_8q�|�1��_V{;�C9�	i���*G�������]c� O2���V��]���?O�&�=/�An���+�ɵ�z2���o��^��Y��I���R)��뭬q��?����������쀏����=W���=�߄G3����ʻ��cѯ?��m��sֹ����;���
�	�����Qq��N����_(����Ea��8�}�d>��}����#3�����&ɔ��4�Ni��z��PQ���+/�/�Vl��GYZrXpLB�{VJ_؁����{g�l�u-Y�ߨ�JƀL�g=��u�Xo�L�9��_j_����\Ȣ�<�~�g,�k?�����e�tK��̆�#I|(u� V�����j�Y����4|��V��ތ��$--�"u�⣫�"�M0��[<��H���X�+��0r0\w'8zl>2�v
򶳄���\P�����s��9��ΒP��>]XݑHSd�ȋ`9��IW��d��	��0y�1�pBu=�)]Q�[����GZ��X�A��I���AUm��ir�+�����q|Ng.�"�q�B�cs��C���� ��\]֞B�r�Q�ee!�p]0I���TR��Cj�0V�TV��D�}WcU����~T� �zUdi F�g��NݹS�Ź������+H;f��K\�g��n���������~�I8��W���bFL��¡�*�#��-�����I��ݿt�>�����{7&Q���V8�QȺ9�LdD�8��x�}-�f}�	
�K�T��V䭁��r��3U���Uw�-'xuRO�sᩆOտ荡Y�z}H�Ƶ6��I���������؄��
'�J��������g����;�z���2���.���}J{$${:��-"dԃ>�5��>�R�����F;���R_\�4����ue�x=��}6Mޯ�r���Il-N'�gEjt��֍<��8}f�@���U'��Ȱ�%!#IP���SKS��B�~���ko���B�C������R�a��ܵhs_f1�}m�6T�!�Rx�b/�K��8�w��l<��{�G���L��	��C�ǡ�g'�����K���B�E|r*��kƔ��t|�gݘM�]�qâM��p]+���~���ߨ���}�A�(�������#@{�"F�E2���g��ٶ49Z?���SG�~���$`����.����;;�_bJ�;=:3��j}z��3j;�[�-�`=���`���u���~1	�Z}[s���x5����?"�1���Ѧ����/b�߱8k��P����*Q�~EFo\��yjc�&��H�^���tn��Q�h���H_5����*�]1��?�'�+'�V�5eI��8��cz�oa��mؤi�5�	�=������ W$U��p�#XT#�C%I8���k�>aU��z�]
t���(�%�e��K� ���~�&$YO97��$s�*Wn�����M��oF�?��h�}5,5%󛻨�z�BP�ŀ���Aø�hK��+���2Vl��>��G��rd�����I�X1/ ��Q'�ﵿo�#ql�g�HXt0(o���>�	���F�Q{KF�uD('&̮/\Ʊ�G�a���Dұ#�0�+3".eG���O�q��Z���q�	��� �������[5@yӝX���3ζ���YIז�+f�ӭ�Xf�=���T�Y���ڐ�\���^to�v�ٔ"k�Lv�T#Ч�n�/�V�ݜ���w�L��k��1�Y��}[ Pz�0�u�Jh�4N	��}����/_ݘ�H��\��/Xjc��	�^��l�P�
�x��Q��>�<�������a��˷6�3�ew8Ů_S�\%O����H
B�̭������HE�$�ۅ���FN=�_��yU�4K�Jtf���P5�?�m�Ϸ�B��R���;��^-�:|�>3�]G��"����.^%��۽I-z\7g��k��p&k�ށ��!(=���yW�1��^�-�x��9����������W$\�O��-����}�\Hjp�y�`�f�7��Τ+K��*6a=qk�(��9F7�/ �p��D����ў�G�u��c) �b��\�_{7�g�e�܉K'�X%��@d�A�L%�G�U@��8�%�wi��Z9��hۉ�����{=f���.j������L�;�ַ�s�AZ�&�e�KR���N�e1�2 Ƒ��D�34�_�+��ʎf/[��[�P���y_�űp�7�rD�Y�/(�aa��P`W�3�V8�~?��j�y���V�`/��V��>ɑd9-�L�sM��lei/[7���I[*n�Vs��-�r�V]�I���8�	O�����	��l:�Z������魙u8����tq�pV;�sHqY�-�Q�
��R��Y*�S�T����>C�Zav�1���"b���t����>�IH4=kMݴcO� �ץ��Ѷ��hs
�B��=N�,�o ����<�<Rro�1G��1^&�$��
�?f �ⲁ����R��mG���B��i�D;��E�D�3�kU�A��K烫�g�3H�(����Z�����=�5���0�B��J�Y��t��Z���gI�YZAb2����XlxVHYEB    4f62     b50u0Ÿ={�RG*�3��C�%�	��o�x썇����ċ�{z6�Q�>���}{�y�Y�E�_�&�#}]Uf -�5�f��S݊Oph0/MS�`�zaW&gch!�W��e*��պ�����js���Q����L�2��b;C\ e}����<���	�( �;xd��hGV��welG���S�O�>Rpv3��s�JaS<]'�j�-ǘ�w�rН]JxƥZ���."}_�{'�{d��n��B����sO�����t�BC�OќU���@�.!���W��U�����fA���*�;�'e�.B���f(S��9�~��xR��\ŉz~��NO+��O�bIӿT��DUE�VT����`���@q��"�|�j~�\_�5<�u�18�U��&�O�ߪD�b�	�bU��g<��DϘ�\����Q��/oP������̛En��*��F�D�U���w���r����Q�Ixg.�+0�O����c���;�a��%ˡϹ8�G�yh�Z����шV�d�f�k�3+|�b2Ĝlz�5� �q�ýɵ�j;��I���5ǬA5����8�P��7E�B.,��.�s�0�Y�=́Ex.�o��)P���r}�g0���zG���,�.1�,��`���6eY���S����P�����=�b�7+�B��q�%��wY���MR�}�{�w~�j`�����.Vۍ��8Z���������Mi+�eF�z��� ����$N^y��A�HYx��>G�~��N��u��|H�A�ƍ���oݼT�-���Yo��Kw�@C}Pو�v��։ܔ����P�$j鮂#7V�t��݋ˌ4�2YM6Y8�h=-�T>\3s7?>Z��,���\��:*k��'�G=�3�]Z�.9�+���D�6Es?oƵۇb�{�<�3��塩�")ر�>ǲ���^'�̖�|�F�����om�Iv����L�au�
����R�wH��H�;p�$va�IdŇ��o��l��i{1����,���{��kL����O���Q���%�Z��W�C����j%y��Y��������ˤPz���r�ԩ�� З�	�bP^��i�|�Q��Ӵ}-�e������6|�¶��B}��&o'!�UA5�S����������S";�˗^��ֆ�Z^����S��"�I
�O�NY��tQ�c�􂲷��X�;�[_�֬�2���l���?�@�r�QNO;r3�����=�a)���T(����+~�	B�J3�յ9y��aU���`Y~����� �Q�R�,GZ S�q��}�|����	C���{��"qP�lc�����)|
^m�k.��i�5��iT�P{�}ՙ�ꭀ��>�����������OV�JJ������O��?����N���s����ء��O^�%>e$*�R�y�n���X�ji.%,��p��%����0щ(�T*a.�|:�7a6���-c7��,[T+x��e\g�����]ʨm�ߤ��KE��ڔE3f�^��*V��DS��_=�ij�J��Gא��d]>м~?�>d�?�*�4�T-�X��pY�~�4⻎G�&��u�k����_@~8��Hb��� !6��a��]B�3�h���Q���������-�.�퀍��v|k�u�	(a<T�:�C
u͡��^4�����q��c�6q~��1|E74���j�@ψa"��B'�w��nח�X
R��4vR�#�xL� � �_�Uo����Dk؄ x����8�6�����OZ��."� ��9���l+�_
R���<r��Eӣ����o�ݙ�#=X��<pB��z�\��a��# ��BbD�3��S�Y�wI��w��pނ��@w��LB�v���������പ54��M՗���Y�N�M������G��b��O1��1�;�N���X�T�ҁ�>�`�'�|J��҆ی����6�euH�Əd��vz�3f�g�xP������}�S�����O�Bx���?5"R��FG�Å�&�O�������F��U�d`zB�-Y]�T��_&b\T�G�aҙ�ا�Tm&����;�MT8�/Q�C�	j�{yG�ȹ������>��[�~e)�io���֛�w��hLC𕕏�V�7�zi��Z:�� �yLL�I�~ϊ5�r������g�U�!$����$���"*�:��==';�|q�@<�KIz�4��+B�UC[e���� ���A��������`P�6�]{�֢�<��/�O�g�Q� ݑ�0I,�|�R��i�z���v�XB���A��2߫�����<�CcBe��	��`B3��~��	���~�u0���ބ5%��ZR�� �"��������� �J���\<�~�0�˞���#��b�#��s`2�#����k���4��^gZf&�n����x
|�����%GB�5�i�P�)i�yct�`
���#ʶ��Axdǀ��ņ�6�G)3��ki��}���h�	s���|���[�&�G��Jsdy�H��ۃ��7�� �\S9�ښ��g���/a�%T�Y�D�h�\K������LZ]Q��v
*�=�c���������j�h.)1�������]c�θ"�J��6�I���&g��'�@E�+�o�wk�kw�N5��$Fۇ5����{�Tf ؚ�`[,lyU22���3�����*"�Kwb��@|%X��������Q�&������og �v�^[1$d��B�}G�M�D�ӄ�e�>q���8y��ƲO�����Z����B�@�Oݟ�:�.!��庮�N�x���垪E)�|�'א�~��:���%