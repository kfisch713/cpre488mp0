XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1�n�����z_�iU�w��nw���q	a�J�2�B \v�r�KA�u����ƒ����e�E�sܘ�3q�c���<��V�Dz��V��������*��0��mc	,��j9k�P`,U�H�nb8L�2)Q a��oqJů����f��Z�fkm��F_�.����7�R_���� o5�剜KUnx�D���u�ѫx�_#P��E�g&���=�5���:�젿P�� )��z��Ũ��E8�8��y�,��NOcv�Q��6��kayn!���r���������gr�ͱ����;��(m���ֳ�2yS^2_hFu
)��r`o�6���?�ᰶp�}sz���FmZ��Si�I���yY���1V�|֕��%3RJG��`�`���?&�6r㣀 ��� �U�A`;���9�(1SP�[�����4�RO{IYR����M�X��GAhz#-\����i�3C�u�C�G��e�4]2Z���G�\^�M��<%h~����(��U̓,��)��p[H��Kf�U�j�7�(�<_k\}*�n��0�^�R U����k�I�[�{�wI矸�v���*/��):���w�Ȱe�*"�#�J��G�i�Yw�����x��ť#vVU(�]���O��1���0�+<H2g���F
����7��0|Q�1s�N�+|�k�<�:�mf�e�\���<���m[���	R80x>��)�D�^"]��ȱ��Dc(��^0�.�^�eR�zhwlE4� \����pF[�$Qמ��XlxVHYEB    dd8f    2160*���Uf�ᄽ��Pn韭Ҷ�Ԯ3���i��,6�hȑG�;	*=?<A�W��2ۈ\A��mƋ\c���#ݦ�;��yM�q��t����pQ��>���꡻�P���K�0�m^�+6#��p@�$|ܻ*y~;���:�-���do+G1��Z�GT�U&Z��e}QI,!S�#�F9>�=�=�;Tm���`W�Aݒ���
�/������t�������$nO�]��0H�T�Y�3V��N�  mv��[�Q�HaQ�%���M6�~���d���0"��)�.�l��������ϧ���&B֟S$΋�Rn)^LN[Z&�E��]�8|_�ʋ�Ш	.��̙�X!�VU�0�r�.��O�����=[�����ɺydQZ�X�l�ॉah>x��FD�L�E�������$�j��M��P�-��̼g�Y��+3�ǜ�i�[��c~���SǇ����рi��N9|��8L^Đn�L7<�~��<�B�#\��B>�&������E�,j0�Q�R>�.�9-�1NV�9 |y���S��賃x�Z�95[6�sZ��O|��F���@�48�)�@�R|b�f��M5g�-0�ZET<BdC��&T�9R$ɋ ��J�Q��������x�T�Y� �*(=,��������E�^���1��Dwf,��+�����Z��29�Kd����� lG@�7qGK%�3�Led#C���?ƻiK#��0&b>��G����o:���ˤomɨ�O����xwd���v`��\�Jr%e�V���v�?���
��!�tY��R�E���E?:�/Rߋ<�4��{z�C�u��97Z��uW�e��m�Aٷ�6�_MtO"�MRA�B���������hj�̱�[
��\���`g���}�7%������a�p}��3�O'��Y�^>A6�!����C��������#�JHG�/�t ڼ�\�?�>$����{�Z�������z9�=Y�����G��
�6�Xfp\go�Љ����p1w���XP��� ���U🛔�q����rQ���A��r�i������,*B�:C|ӄ�$��t�e}���S|D�&4�p�45F~S(O�uD��w�(|�t&��R+���r��<��w',_�^�cE:�bh'?L��{,���T��i���\b��U��b�=T�A�9F1Mn�i�Hz�hw��
'	����
��[S��s��e�ů�/�����y{����waC`d�r���="��|�k/��l2�j���
Ԯ,a��6�7���(j���V������RU�����ϼ=Ve6 ��QGhО{D�0tn�%8����t��������AYY�{�E��Q"#Bb�8��b����>�E����-���y��2DA���91ID���~�N��]}�ۓ�j$we�a���Ɋ�Fᛀ�r���2��Ш>^�-�j�ey!�O��Dn��<���e�@*㿂f4z*Lхx�S��0���H����������@Ŭa�._��̽Bx����Ƀ�;���i˒Y��Sꭘ U�� �S]tw�XiI��qz�&�#֚2k��yl�]�%��]�+G����g��@x���/Z�q5Zo%[��2��@� >ۦ"8z���wЩ�KL*s�S#�q���`10X�\J�6�,zM�Q"D���x9=��ik���\C�JFͥ�����
�e�w ����4�cX;H��^��$חLN�Q��0�)*�� ���<��/��tFx?	U�;0�o;_��l2H�3vjf�1�t��p���c-��e��U�Ju��]|e[��#F��q�{�q�A����f�(�����b�m���G��a�z�sI7nm�:�� �����B�O�']��ъ������Nʥ; �o�/De���x�maH��&��^��F��I�`��Ac�|�	�*����E�{6l߇8��7��
��l�<'�s����fF�{�S�Q��1�#�2\�@��u{K�ڢ���l���Nh�?�ͨ��X+
��HX�y�K�d�?^T��SD��(SiV�,�{l�)Xt���DJ��{Z�,�v��#5g!	���1!�OTщ�O�3-�����Q��>Qq����R�Ʊ�i�A�[�;�`��B$O���^��SN3����;���r�H�p�N��.U�^o��/Ni�a`E��9G�u�5>��S.�ѹ��?�=�,w�Pl^E�aT,ʔ_�A.<���u��
��{8���_0�O�h%�]�]?ip��$6/��>�I�拺$��yG��h��m6dA�|��.��o /J�����ٳJjSS��Nn�@I�W��@MǢ_�h�I�$�JF�J�_׉& ��RIX1W}j�s� ������]Y�8:�}�$5�����v�1`�k���(P�5��M�p���!���׼��� ��OV-�cM�M�V�q[WI� �Alee�~��R��[#-쇦��E�?����n����4�%�c�� ��o�xR�5qjl���A�A�aK��C�������M�Y�>�����v�j�'��������>uH'��G�?Y��ߵ�k���藶�u�pj�*�h�j����hi�}5� �l��� �ײĎ�����V��(��>f��\0~N���6�P��� d""�\21�E��{T+�-B �ꮁ�w~kQ���(Oo��G�+`�Zm}��!{�9�kכ�V��=O���s�Љ~�	o>��]ޞ����x�gB��˃z�Ţ��g4�T�/�!���m'���CA�Md-B�]�Ӝxx�sV>��z"�?��X�"��Q#�*�A#�����D*	ta��b�=�? ]R��k�H�D������{��x��m{���FE� B�}��WC+U�uǉ�Rj�L����-��M �	�aUè���Ub}���T 3�J��c��mmml;W�wb���Ws�O.t(�'�6n�Ȩ��t~��Ӵ�cS(ڻf�c蜣+Kt�ʏ�|pj���T���,Yǁ���4V�@ِ�|l��Z_����NJE=ɕ!�rެ�V�P���ǑFJzA�t�
�k�����E�b����i���b�0�:���8��ܦ���K��A���Z�r|�f���v�����|�����Ugif]E�_��Z^��N�
�E����Dzv)��d�)s��*kQ/}JÙN%�U�e��ܹ�xIcx�޴�d'�<C�w��q�D�Ȏ�+�%
)�,�=�j���Ie�Y��z;(��'�ȺZ�oqq?������C�^���-����_���S��(-ә�"W l�]�aPK�T.�� �65]�o�i��������)�P6������s�E#-P"�P��I�]�#!c����ב}��4���E����]��I}�y�t��ɞ�@��a�}ٙV5"M&G��@�	�.�����[�y$o�!l`��>�j�A^1{���K���2Jz��%��]q��:��Y�st�+ÅǞ����]/�fU�
IY�"��m�{�G�̫��"�׳�=��v	v���
�D�#�K;��F6&;�/���v���\>�����V�-�5��g#`s������p"� �9�\�F׎wx��F~X�Vd�Ƶ�R=Uf�ޮ�
�^�MG�CQU��t��ܦ��;�^��y�����e�/B��N7M
A�>�(q˱P�a.�eНP��j�HFb]�&�u5�T����M��h-[�*�,��+B�h�h��[?^`$R�u\��)2��b�dH�:jA��&a���/��դ!�T�J�Um���3���pP,$�/���<O�E�"�I�� 7�c9*�,�N�!�\�[1켪�v%ٳ8�sJx0r����;�eByLhޓЯ��e܀�����1�p��T]�1���x�h}����� 
7���e���r�L�a��9_���h$A^5EZ���U/]3���qX�l0�%F�Q.�+���[q�T��$%��3o�?��@7!���RU�$hYHu*��(}�KkT���.�"Ѝx�*���l#�L2j��%��S��������Ɖm�^#���E��E��)tp��`	�]��]y`�|�C��`�M��YY#��ֲM�~�@kd�QG!���i��7v�$��l�� twh�NC�����6��T/aQ�j'J�,f�N��dG��	wư8d��C�LR���0mƟ�z�A1*�)e�Q]�����']���4�,�8�[ae�,{��(�4d�Q��i��.��"(n��#� ����Ҙ*u��ޢȐ�\^�����x9��M�`�ܳE.�N�F�ד��������_���p�����b��Y���L��51A���cW�g��i�	6�F߰���>ǌ6�	��,r��̋/����rK�j��@
�w؎�	�3�-&sڍΘ����µ*Q)� 7����y���/ٲs ֻ��!^�a��m�Qę��kK���Oz�~�Ǆ+KX���=���8*41�S����������)Z_����u���i` �_�7��kS(��T*pa~≛�9���օ��<-�Wi���8�����e���0Mo(��VRa�b(�C�j�#+
��6��H�t�'��>�3����S��l�J<�/W�-�R-h}	� �J=;��l[�~��FI_���Cyj䬚���R�{ك���b�h�B ���oP%����9"��Yӧ�6�VPްq�`	:O�>k��CeT�B� d�,�*U�1�D[˛��؝���n��д����iܯ�*]v�4�n�y�y�u�-�H����wk|u�.���1��C����c���k�%�l�!^��";1X?2�U�8h�:����9����6fY���2߯���0
A�L(�V��������L��&����� N" ��*��v|M/�e�u�e�;�b���H�'@/~�|~͙��N�A��������T�^���z��A�m��A�0� dM�o��D�Ub�u>��:�V�������D���l�'� �VZ���w�+��]���S{屙�}4�����$Ld�O�Y��f:�R+�S����CK��1�"�ànF?�%���Mu���?o/�ECfJ%�Sk]y<�p���'$��c�gѵ��d�~�<~>�a��b-i~ꞛ�/7�=	i��x�v�MAw�4D����Gl�wRj#=��r��h?�f4���8#��+R��q��ZL��C��x����3�XcY|`Y�H9Is�dt_ ^���1���Yĸ������-�똵��ޖY�8e�����Z�Νo�M.5�""G�0)ϵ���;5��`���*3�ᙫG"��%d�=E�D}4ɑf,Y�?��"�&`�W��4?E��j*���_���G�}�S| ����L��zj��%+���{� �#�}�I��v~[�߉bn=�$pP��.�̡M�O�'��&�#��+�&k=�6肁֥�����u��b�Q���ͷ��3DCF>�b;�O�6���K�:�����G��2W��44�="/�.1p��U9��
�o�u2�\Yj}��ӣ�u��8l;F��#�:5R�P�Z���x*)H��QF��@4ж���z�z�$mB�HF�U���o\t0��mv������LH������͟���L�"YKyH��U�;��T������H�N���7\%Lf�΁���@�Lf�ڒ�`��O�[%�e;0�ίHH��à���v��#��ٌ�^i^��&��W����K}�4m���b���Ǐm쟞ʝs��"��^�DJ�����C��xKw�:W�@y�}�=F���
��ǑGّ����PB�ezT�>�Z��,!��
F���p��H��	U�߭��t]2O���D���.lA��.�(�{Y>���C)�f�}B��!d"������6���T'�NR�^�c�{$���V!�3|�6�`;<uԩ�O��-c��T+�j%���}�0<%�����ݢ{��������|f���'r	|��_��p�Q5ܦ-^=�8V�I�A�c�������ɱno(C�3��=y�	��nKQ�������y�1/Xf$?��B�������{�C�gKMy�t�G$9��s�$�N����C������y"�^+ͤ;q�[��m�.R�8��+�G�8��'^X��2-��D�S��\5�^�our'������u�o�u����#������ׅ���z�6��kȀ4�s�9!@����)������-��o;��4d�6�������H�!u�L�Ά-=�>U����xxYy���\���t����:���8-�c��UKe��PVCL=O�.��[vz�Ht�^y����������nP�������pr��e�(^�<ևC�����g^q��=���$������h������3)�Р�a�2�};z�''{Y��Z6F�u��Ծꑸ�ACm]^��5]�ӻ����-s�^��8�Z�����L�T<'7�u#�b���F�m��d�k��&u��B��o���Z�p����B'�-[ ����M��AGŊt?y�}��"ϩc�2����(�\�P���!�S�"��6/����C��V^3!�*��{}�+��!�#�a%\�+�k�Ubȏ���C�Q$��-m��<���u�H҈6l-�w�Xk�3�}�PF����~њ�Jm�3�>��G�N9�7k�0Al�u����з_ǇVg[N�{4�x�f磩�Tժ"��$�R���ٴ�0LЪ��|��:o��C1��T��������r{9��*�NJ4L�s��zLFc��j�5!���:���Y��@�HW��R���+L�`d���ק��Q�#y��Lo�ȟ[��/5���#{��ѶP�������k� g� R�@�	��v	
���������o��Ĉ�*�;�95�� ,�􉆧��2��m��B�+��a6�N��"
�
9����k �Lk���T�`hA(� �A�\D��dg��Z�S�eH�T�g�X���c�y ��/�ŅR����tޅϏ�]��"E�ܣK���++#��>t�?���f&~ ���ը�%�l����/�L�A�z>����ܺ��ŏ����g��1�d����c*?{��uEA)¬�w-��� �8��E�5׍���$S��'�
��j������ηHDJ��#R�L�:�Q �����@���tz^�z6��8Q@�f0�f��(?b6�ź�Q֯o8om���Z+�%�0Cݙ�ߗ%M �5�D�7D1堍H�ߦ�������-Νsͧk��P��b�?�6\�v��i.�p���P�8��&�gEM1������ÞB�Ǐ��*[1�7Eb@x_���*XFe�Hj��˜0��6�
e��Y ��|�p;���0��)Lr����}�Z�"x��	 ������%�z��vy�>%����5R�´����{I.�'�)Un�~T̟IO��/8u�48�ҷ ��Ր����}��?|L��������yjO �x��jDGػ~jJ�e�o����X3�������`�i�lL�����on}�Y�a3ܲ4߲�oV@+tZ�$@V/�i4(��v'(�7��q�|�͋�;�Af��&;�ʀfi�@v���������fy� ޯ|�֌h���
�͏��Gy����O��/D-����~Ly�-\$�֎/��-�?�1��`�@�r�Z�_�)��J����Ë���!)�@�R��(!���~�U�'���zZH_]��+����2���(��q�y2���x��|�I#L��Qwm��E��%=���wn�t����;Gz&(��89��{jC&*���о!���^} �{z\%���u�Ĭ��̰�q�GW$����X�D�����s�5����SB;a��@��ٶ�W߇��Xz�Q7�������ޮ�o�Q~$�!S��n��Ǿ��R�;��
"�$�i�"�6�8:�h1�Gj�+,;�������4i��J0Ł ��(Y:�A�R����1i�5d6^��M�w�,�&�Vf��ʦڻ֋�IWcL�����HX{C{�XH'��iڒ�U~RB�5��N��%���ů�,�]@���d0P��y���`�8�(xek�I����C�C*���h�z��=sSݭ�����f�@9�T_�2ܖ�kpAVg�*3r�&��L��b��3�Ӵ���zݥ_��������z�s�	�گ*��+5�A��*���C�m��E��}y(FcGT \�U>/���!MQMN�`ꩫ�֘`���G��.�����J�>�F�����Jl�	�a@�Դ��&+:v= T����I�=\�Z��E6�'ϛ�a��p�щ�����U