XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���k������~��q�`N!/?�v>��-R�>�l[\��,A�+�r@ĥk����ə=K١G�MP�\	^S���0����7sFᶪ� [�Fԏ,�v4�q���Ĵm^qv�6�����$�xcS� w�~+Υ�\�~q����1E��q�{Y4��5��t�
���q�/��\��ّ��BX$^�Z�y�}��d��
�Gv��XqA>���F4u��R�G�xo�V���/ ���͠��tBs&"���Ʃ�j��/^یW�4먩�B_�q��nŶ'�Fp��:>{��g���n�^�����(��x���V.wVd��<H��7�,�/�m�����!�	:�$�p>^�*ԇ�W�����>t��y;\l�v���1�FM��xVrZи������0yw��C����	w�|D��������Y}�B����D:���u���>|���FzbW�S��=v%�x\kc�홇��\���N���!zI%�b-M��h��z۲�	.�`�� ��u�݈�H����p*_��0:?b�S��jӢ>��C���� 44�4!�cp�,��1�ZGCT|/=�����o�u����X~�������,1���I�+�soJ��Au���R��Q��G#~�Ԫ���1*�͕F�b!ŀ��jq�i��.�&x�2�
d��lT�̖����������	�O~<	�jL����x��wG�ڊ�c�sb�j��a�TrZ�p$�������ɯ%���Bݥ*=���2K�j==6XΏ�s��>-XlxVHYEB    fa00    2040��O���/��'���_��ꩊ�OA.�-��x�N�#�C4����+Q)�	��jLE]j�|jZ�G.���� s���(i-L��r�s��r��P2:����$q�魼�1�Ϸz��L�:g�J��T�Du�nG\E�-Q�u��?G�J�^d}����r;6��[��2��1�;K%�ö)�]$	���nd��(�zS�JV�Y!L�eJA�iwuE���u���	�������3�F� #����6a4��*��h�b�r
�M�ͬ�g�:B �̛�-|4) �&d���%����mT�0�E��{��7`W��u��A�7�۩ͽ��'�W�zBn=l=�H�4��AZ�D���d����Գ��.G`3t<Z�`r^�I�j��#
^g��?E�x�J��?yR;����Ka����)�A����-���A���fQe�v$O�Cߏ^/nള��nya�-�"���@�v���l�.�C'�`�W�L��L���]��=BH]�p�F\�Q��3�^�B��t���s�"��o�mytxJ���E>�6������γt8�H�C��q�oj�*�N�P������-�.�Az��S�� &T��z�"Yc���5��$׫­�����0���X�X1af��ɒ�@ȶL�PO��c!��9��	z'�~k�]J���yaC���Ϩ\pN���i���G�7����!�Z��s��z����{��sp|���?aW6ǫ�!�%)Qfn��2�g�g�q/�XX8�P��6��k�,'�ψ8�fw�VF��@���4�'�����wP�
 j��n�5ݜؠc����W���7��Rus�#���p
 �Q��{V -�ye�����rI��Dh� �ᄷ�qp2ʌn�	��"a�bϼ�/����9d)b�2T`��U[�
�?�ɍww��q\$�t�l�򱺭�MW^��?d��I/��L��z�W��&��λSW��c�'Ng�;{�׿g�Rg�������[LP�2�C���� %de�Y���2`�O�c�+@��tT�KKU��>�gfb�Ȳ:�&f@�k"Eq�h�%"�:�`��n����	���g�r��K�ZH���nVG5���"U�.׷�W�"���M�����6{��좠TBGЭ�N�䷓k���z'�lzl디aQP.�����z����̥�}�u�5�|�4Z��ѧ�V`.�Gx�Ug�����Uր
�1��A��C@����	�����wdP�v�~����ۍ`���Kd֌)C�U����,d��4;^=xΫ��6;Zz���>����g�Q�l~�>Ն<g9ep��_������f��\�c�>-�=8b�	0���Au{#��y� v',���*~�9EW�v�>zO�T�?zsB|��E��}͵2��x�g��E��k��.n𘠫��=<Ա�rb5�0K�m�O�B�ؾ���ӿ�:��_3���	,�u
���	P�͗W���\;x�����ty�,v_	�4]��#(�b��>� ���ڏwM�����<����^��G2��D=�\��(Da[�g}�ڳO@Ŭf>�eET1~�=ZA�m�9�C�cMQ����U9��G��Jo���M�Mۭ.�,�?$Mٽ���PN��77I�)���m����վ�HPZ�G��e�#HF����!-lF��m	���������J���B���ieH.ߴF=���l)v�!��`\��V����ږ�^����|�����`�.*��X=�	���>O CY*a���;�"*�B�ݢ�ߤHw�Y	5�w��v'C[z���.fo�ɖ1��_{�D�&In�w��%J��)~����9�Z���6p�w�[�C0��|�Y�Q1�
AL7^)v���	�u��*��~�B1�,�� iF��i����J�QP��>᎐�:܇��U�0c�+��E֮�m�$�%Epy�M�N��ҿ�ty�د򫍙Ȇv�&ظ�6��i�\>na+"�����8����
�Z�؝ˎ��n��p[� ��e�ĝq4;	P��ϒ֠Cʖȋ0xm��Z�[٪ h������$�Z���t;j��o4���X
B�Vu����n#�^  �k�P��4���`��gw���InQ�k������9·X"��h���8��}�uKP#w�{� ���3>$C�b}*��ׇ��)�����Y�P,�(^�.#��+ 	N9����}��4Pn�'^�m�3��lC.�C��v�ˍ��p��H֖���/���Ķ�c:�%�J�'$R.��5���ձD�X�^���Sz�X�רU�裀�c9�1`i1'�+���>*�-�I�g�������fo�" -�+�A� +#�:Eu�T�a!='����h�x�#����U���"_Q?�[& P+'x�S��Z*��A���X=2�;�'��`|�`��A^手��Qp��҇���g�uu�m|���a���3�p�R=x�{�OK�<���HA��aQ��ׅ��,D^/q�]��>�K���W ��#|�w�+�^.Lu1����m$��i�_g2'������d�*^��9,���wf�;�G�}��T���*z"���Pֳ�h��g-W��TU���ð�*��6�����\R�_T�r�jA~���/+�L��#�	��Ax)d�:���a@<۰�V��{�(\g��s�C��v�s�^9�FS�h�������;�=)X�٪�����b,��*�V( m�@�b -�t=��u0i��!�@y6Q.��G��Ia��]J���5���UA�N������auB�u81n��2ef���@�SY&�l��^�+�������=gt,���)���7ϗ���!�;�|(���V��󛶰�.N�K�S@�cޒ�
�_���W{D�\ܢb���ԍ�,,��?N�7�=
�S80ֲM��
5�y�`���L���֜��׿ ��3�nV�Uȍ<��r1&�PB�,�)Q�;�)�ُu�d���4a>������ ��1��a�& G�nJ���Q�D����Y���"74.(��B81� I��>��+���1����Go����|]����ǈ0��y?ʂ�����.zV�h�}Kk�J��kY�����,��?iF6*��P���RO���ҽ�k(Z�G�B颩��c����N����)��i�b��V[?N�yݕpP���=�������5���
'F����Q5|�Me��HB��ʁ����߄>7m���_�b5��������y,�j�B<�2]Wuq�-r{v����D9��os9�t!l�,|��E�[���&,姭d�<���n�#^��3�$%�Ѐ�������%�"�*��l�@d	A�r
�l0����쩬����6w��_I���j� �׶�=	�݋�F���@�,E�֬�t����ش;=l���-6�~��Ň����~�TD�fWfka���:��q�Ea�4��ۤ����9JBl�����.M��ї�S��\�A)�`�O��� {9�]�s7���qގXF(/�_�.������
�M��A��7◵ĻO�Þ�X#� ִF����w�M>��\[
i0[�~�0�4y�f�V;��D���ZRּ*�^]-�lS�H��c�3��|��'� �lQ��l��#���;(��P����D���A𔦮<qsM��I.�*��5����sA�'�]�\���a�m���vO��9	���{� ��~l$���.7+������b.�H�Ьcr�9G�@����ǥb=V�O')[�eK��=q=���<�1S�u�Q����\s܄"z��t1�َZP��n���U���u�s6zC1�r�䤪�z��\P��\n#�HH~����RTO�JC�}df,$��;���Uѐ+�-��� a!ڶ~�ux�ةM��y����D�o�Ld@��ٲB:�嫖"jI�O��4���
��0��e��u�5��r_�Q����Ñ�����.3nOqvG��f�,i��%?k�J��s�!E�Z�X�����l&fД3.v�r�< srj?��m m_��S�3'E4�\�f!.�oC���>w`ʽ>Qj:�+�5�\`��ܶ�پ}4�:��.��Y��i��ٓ�q�oW�?�A�K�V㎮B�Ϋ���/�~(�W��~��<�R�;ͼ�i�D��E��c֖Q^�����X�h�u%]ך�>}x�!�c��b�OD�f��z'[�c���\
�Vh�1������c|#��L����U���0���>5��~�X��Ļ� ^��NQ�徙��LUV�P��24�j�@���*ueg4N5O�o0�.N)�z� (1nP�OX	3�7���p��gɗ���^>:��:�6�(�H�X<^ 9�ڨ��tӛ��t�Na4��!!UN覉�����\ ~���.v5����W�|�6'\.��ċ��[jgA��xdlo��o�=����KMKN~���(���@<���hat��l:Hz�I�ap<�I�soMjGW��-P�k��{�ӕ2��:�ZuCÂī-9���@�
t��$k�?r�á�:��R�uӔI�Y�)��yM�'d[�m.QPG��&wQ�͚)&�bCw�U�"�Ħ�[T[���0!�h������p4�Q��>@��Dڙ�-5�(�+Q���+�
/��g����Z c�O��q��X����q��s�A�����t�2+���+�ȇ�4�	屃�*����@X��]m��p*�a��N��Gy]�"TG�X�/���:y�.��@s��ǮY�Gs�p��`�(Ƭ�^��2�B
l��L1/�{t�^�����`�bQ�R��izNcap��&QexM�LP}Sҝ���{*/ ^��$�4�R$X,Q�j�Xxْ����5���[;�pW��%���9cZ����#{�_��DM�����J��¿���a�@��Cf�C�ȝLf6���"�j
����ό��H ��ߪRY%��h2��đ_��`�b�\N@�f� ��,mЛ�\�Ka�Sp�����]|e�ݎ��j7��M�؊s6�x�=�k	p
����c}��
�(��������k���zq�~3Ҟ��-���N)7Ƚ	}�ҟ˄i�H/���G(im��h!��ܐ��\3�Z5��
RkH�]/ l�����O��*`�2Po����Q�Mog5��h��j��]}��oѼ,��u!�=�g	�{y!�4��u���C��~�9H�#t��	���*W��5;Cq"��x����RQ"�L�+�	eq��#u�o~�7i�NzA����:�v!����w�}$"F���`�$"\�P�9��꺦�������xj�j*�1Oދ�ڲԃ�aV1>��kB��R��Q2p��{w{�*3�|��l�@���8��2��U���f�HRЋ���7��֤����pR]����!���J��I�*�G��YǼ�D}��8GC� yZ��}�.�q�����W!b��eL�,x"3�G�>U"��HnX����:�5�'����Ȟ�e?��]C|����x�,�ӭ�9&G�
[��B���X��5b�!o���!�Dt�9Qy'�F��C�6�0v��k��Q�~�ղ���W���4�ʹ�@g��+�r�Ӊ3|�"�[%��~�
�Aƨ�b�����x����W�|�[�7���ILA�|E�,%�Os,A�gJ�x����z��,O���	�`DB��b�ŧ��E�M:�����#�b���F�Bk����Rn��&���N@��̴� ���}�3���=^�u���1�[m���]d�gk�|h.��#E�<?�Q�=�y�_�0?�@�i�]C� 1w��'���T���Mٰ�xu,@�|����WM~�mKɊ#��G���՟�����P��r�h�{kWӳc�-hB��#W�fU�AsY9�uxB[-��y�]�YGQh��cɫA�s_\z���"�Vq��Y��-��n�:�ш�z��ݶ#����Ae(3S��}�IRJ�=m�w����#�BS+=�5eBy`te�O!�+(DF��s�/S�>E���Cr9��Hʊ��F&O�|ч/��Y��֐�G6<�J g47R�S�ڌ&b�BrYb����@��h�,���6������~q��O����6�쬽��.�P��V��e�Ҽ��9�����(),��3��g��-�#ҾDv�~�'��@����酓O���g��(��Q�`�����Ac�X�����q��̤.(̯3�>��n���Uǐ��t]��.F-b���º�"c��E
��&Wt�8�Z�(�C ��~ΠFgXUr�o�%Ӓ�Hk.h�@�}$p�;LӯX��Q�4���U�1� �7�i��:p����~�xl
�����%�f���.̼m��8��8_�w�p�K郉y�o�*h��kBN R�<�����:�Z	d�'����}b�:�F�o^8�ȩ0��n�V��Ln*���ϋE:%�01pT,c>���a�哐Z(ϥs�r!N����,+�v/6�g��5����6�&ћ%���M�Ӏ�����uHf�<
&<�9��B��c�W���ǵ�f=�%�2&^=h��l��٤�DG<z4]E�}�4�Gk������e+��0��Ak�]���\wZ�*���<{0�(gۑ���8�<�:_�Q�v�#�
H\-P�x&�f�w$uB֧s~\�2����>��Ք�C��g�o��|�90�}tꕊ\.���U��H�uM�e�0s�Og�	˴����ێ>�oI�^���D,:��}!��^���b�\���Thu������y����C�4��R��+X�K� ��x0r3E���uE�f��n�D���ת����`<s�<����a`��(�)�����Ј1�F<����?���V@���Ӡ�Z��G��y���ee4�
�=5:�m2~�n_f�=,4~�� 8�;����d�G2�q�d�G�{��[���f��:�JGY[�q�\(���>ESU)ԋ�`���n�$/�J��٣�ü	%��j���(#.&l)��_y������:�	���ַݿ\?�(���>��3CM���¿��8FD8D뾄�C�z,�'�ز�<�ֆ5{��=����bT������KK�Mh���6�\R+��=I����n��
����p=��&���sLOdi�Z{�ݘ���M�����>�s�e�w���te9"<r�ԣ�`{JA����@vhnk�3�2݁*��(f0]&M�cF�'&a�5�D�y���)x�":�PjJ�d)#���ߏ���"fFh482����Z��u �EL��҅\Y�}�F66@<!�W���EN�x5i������to�d��/����3�E�k����A�KߪJ�A�g�^��He$��]�qmL14^�N"�F�!WǊʠs����?!�A �$ɎoҀ���vr�~��u���Cy���)F`��פ%�w�u%u6&R�1T�J#�%���'WP"�5�Ϣ�~��q��A�M|h0^vx�#�zнz�����H��Lb*bhl���c�(\S��@�E�
�Ӻ���/�[�Ȥ�gڈ��(�>�p?Nb���������쵞���(���t	 ��V�����ޏP|W#�Jan�5��a�?iĊ��f/���	�:�+��r&��9�MI�[/3�H�}޽�5G��Xs�>���(�d�ֹr���ڄXo�H�{��؝݉��n�`E���w�qcT�_�!�q��+&��I0�UK�~��:�L�y'd�Mf!�r[S�W���O:'S��\�rb/�t��~O����1%�:�����C��XK�b"���xT���y�(���u���qW�Ƹ6�0����}m�ֈ�E�v�m��e�Χ�VaY�)J~4�wU��$Bgr���U-�)I�z;ꖹFK�3�}|�n���Ӊ���-lG(��paT�:h�*ZG�x%�P_O z�p�p@NrmD}#CQ�v��SJ���3����)���Kz�>g�����<8���E7�.*!�J��5���A'c)'.�aR��1��$�i? ��9��8`k�yEr��xyE�\�TǏ��M�XlxVHYEB    4f62     b50I3"4�d��R�� d��:RdK�B���+ƣ��D����c�L�)ߪ��[�y7�}Jm�#��<����n��c#`�&l?���"��n��Vf-A��&�����^w��2����%�X��1��7�4*D2���`���[d���5~ǆۆ�n�;({ܑT��M�������	L�Ć�|�&s��K��p�9�m9d\t�����q��K�!`~ҙ��������[�kO��Ώ��Cmjx���P������l�I�S ��Yi�b��������u�E��RHseX����Ӌe��N��j��zH�7uHף	�j������7��t���1�w�Dv���.�H�JK:K�c}4i�m���A�5�TşV�����y���+#)-K/ ���Y6"G��u(,�O���}�N��h2���J���)����.aq!J���8C�W�
c�þ�
�l��A�`�Bw����D�#~��t�j��oQU��!DB��$,�^f̺MF*��J)��8��;zf�g��.mOX ��>�`�Jv���3�R���6�Qo�zCbuj�<՜o	k������t��D��8��nFy�'�㭢�-��5��5T�� ����+
Ȏ��JI�^! E�F91Q�/��fhM����lg9͝��4��8e Ԉ��KJ�Ih�|FMf������W���(*�0D泃*i�H���e�����(��)C�5[�i��4�;�C2M9�Ԯ� �7ʳ�G1��F3���m��As���~�' �{n\]�f�U�񪆏8CO��A҅�E :n�3c���AH�a�B�������.�>U`u@:Iz�)S8ᥡ��$2�ȡ��j`�cXE�m���b�B�}� ��Z�^ߒ���Av(-�9����^o֠�U�O�iU�G��+�q�T]�%ImU�����
��;eh���H��%�+�����9f�*� ��<�*~6�;��IVnį��SL��`6�UxXU%PF��c�t�&�(�n����ɷ��|0\�����CG"�=FA�����2���y��D��<�+d=p��������@ ����Ҋ49Cqݣ܅Dh��2&D�Rªp���Ob��Z*m�Xݗ�qt��?L��(���o�5Z$Q�����
k�7mÝ�g�P��:TB/���y�!��&
�M0-ęt�R{,�$�".�Qjz��1K]6�L6��ф=��$Z���wsb��d\>�q�#8��\���&k��ι�i-w�8|Pt(^Py������D�y�O�x�<�����\hI�S���=�:{�v�	���o��k�q�� )�"�?�N���t��Dp�x6nʹ�mL�G*=//�U�6�(,�YA���Ja��ج�k�>�~��j0ߢ�5�����I}�H�B�8����v|�c��ge`<-W3����αH2�/vx��[���x�F���q_��:@@Q�)T*��c�=���Ԇ�$)U�3W��Q1��1~��T=�v3�i��ec���7ク*hJ.R$��`�]����/V�5Pp��}WM�� �b��aB�-�Ŏ���� ����%%��Ա |t��!rSP�UB����l7�<�p6	}">�`��#l
�}��M�1)0��x��^)/eʴ ����b�h��cM�d�H��!xFq���/p�v�PT訤zR(�+D�c�_r���?fP@��g0�$�(LM�����#xCp�
j��|�0!��2Ƞ�W��d�2���.����)2�@��]�P�ؐ+�/����~���S�}�ږ����X�+�j�XP�+�%+� �ۛK�X	&��CVR�o�f�Щ%�D��mx���+��Zp�W9qlz�q�7��Сv��A�����������]�=bIl�9g#�\��\�	��H��~S9��C
 �R�v�L����y�T����:��o�{�1�}/:,�:��i�y���A�v��:ha4-��*�c5���vr�[����@�C����.\��1��v�S1��Yqq������+�z�n��p�/ �@�m��=�*Z��B��F��-x�O�W�>��dp��<��0�z�E�	�PЊ�e�|�ƚ��:%n��]�50)��9��Xi��m~��@�T[�U�W�^��.I��=��h�����_Eg�|)$�Ȯ�h�;Ft��=Z��y��׺x$lto:�±�.K��<�RU��෭�#���v(�I15J�4�y�fG��Ŧ�d�ei����;�w���7L��֣�{;�S�
��]�z�ƈ�������1�+�K��4�F�
�I���}�b���0���sXҤ�{(�{�OM��2���{ �=��@3��=�#�?��ϧ��er�y��΁:��	�u�����w�q�����OZPFJ%���k�n�礀��(�E�ޫ�(+y_�ԭ��r�?�c�B�H �X��G?h�=W�c�8�����ͤ��C�����i�?xaԸ�~��ʹ���+���S�Zu���~b��)�%���NR*��<���C�FL����&磢{$��n�漢�b�9R�h)�|�T}Ԭ!��8k.�6����@����_|��>}�kԼ&hkw�ƻ��?4�i��7Ո�k�|&91J�E��B��M���sof�Oj��Y���'@�ѧѝc\���%jO�}��Kjzx��}���G����ߘ�@V��8E�?/ 7��YQ�  ����7�_���6�#���C�ȷZ! ®�(i�I�^XE٤������(�g��@�5
	��W�B÷H���b
w�+gG�X;��y[����n����>�F�m�l;��b2�g��:�+�#��\		�����