XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��uYQ�m��Ya=��#��t�}��=5ŅQ<ÿJ�m�H�P�Z���V��
6��@��`��=�?��҃�1w�B^���-���v���@L"���u!#�נ�QE������Ԣx!�K�I� ó���M�r�f1����y
�!vD_4~� ��\���s����I7��\���eb��i�4���t��5GR���_�A�\SV@n !�����7O%6����h&�"m1�������
�gTL�w!��3I֊H��:꣫�)i������9��#���Y�aF�1�6�jVe��X�d^
rb?�b8i���vv9AX�g��(
�q^v��1���%��JBW�%��,~�S�Bk�X���k��'P�t�1)��E�(����ƫI�O���@��'ʡR�T:���j��BNz_�WCk*cV9� I�؍�baBd܊L��4o:�ܢ���кX| �cH8S2�H*���^w��w�/$zL������N�@���&w����gUM"��b$S���� �,�)η#"�6�3�)���N�24An_&-r�B�>�u���VԱ�����E�WӮ����y&W�~�K�{�I����@�Ә�I�\�7Or׽gR�[r}��m#`��>�s���߽����d�	I��o�}Y�E@ϛ�g� H�I����D���[͆�W���:VЭt�S�i2,;}�t�D��~l!���{��A���T�N���PsQG�#9�9��oL�ynz��XlxVHYEB    6346    1790l�ώ�2�ґM��W�̺C�K�o�o��
��\��}���""�띱<]ףv4�5�F�[�E�Eb�S���j�k}2m5��m�~��������Ĉ�}���Y�Av�e:E��R�/����G���-O(���÷�U�Syj���ig���	�g��Z[,b�uWZzQ�v*�تP/�Ir�r��l�H�ږ�<�I����j�f�M�n��!�+�C���]�;d%ox��E�}=;=`�[���OIJU����Z��g���|�,��'����)�@�����7����G�M���B�܆_���̤q`�x�`|�49��>�*Q󧅪	E�{>a��Eq��4��l�Qj�`�a���ԁI�pp��U��	��@������<���G�����X۫�O*�Q�9?d���%�vI���LU�og��+*��
&�LS9��ft�ȉf	a��'6@��?�+a���c���)lf�lT�ȖF�6�ڂ�����v�@a֍j��c&s�n���a4(���n�Z _�q���6LM�@��m�'�|��H��.��*��A��Is�b@��m�<��w�\A�6N�m}��P��N~���y��._,/:F6�{o�%��W��`-Xc�@��y��ۮ����
���"��:�ܩ[�$�(km��l�G�-��x&�W���lJ|l;"]5�����_��l�̚���[��h�	ƛ�� ��.�]��$�:�3�Kvxg�H��9^Z!�B��RR�Y�_����-5���� '(9%�hh_�* ��R���g)��j�C0 n[����N� s�4�i�[@=[U��p4�We�ͣ3a��<��`&/��γ���kSn},J�a��`�O@�'�����'��AF#�}�Ą^�J$)�!�� }{Ph�|�:���͘8'���'��X~���Gu�;
[u����\i��i��m� �U�����n�Yz���l_����V��Xu�	p�9]��R#ʺ*(�؃���<�>�7V���B�.'�Rk��g&=)�? -�o�i�¬��̄C��l�*�@ޖ�l�+��
���]��R�Z	P֔!��POJ�Y�2�T.�qc��J�qd_��wS���E�Ǻx.[\A���H��uH�kG�+QM��W���{���Y/h�����T��������yY�Kc���Օm�N�I0y��
��/Do=%[HFs�� �Ǎkx)��JE[����]K��c�:h�Q7'JȒ3z�/ @A����۩���K#ø&�ų�l���~yQ�g*�7����M��^����u�����}�擀�-�L�8U�_���U�O( (�@Tf)��gHfsm���W�������o�]\x�$�=��D+m׷�c~�#~ԑ���������%���l�r��!�n��:���V�*{P��G:��ٯ� n(�A�c����W�_�p*㋩�/����� �9o��o���]� �q�9h�
O���{��做�X�bݚB=�t�N7�	ڰ��B��4£���q��Z5�V�A�]��YA��-��$�f'��k���g���w.�����ʑ���v7��a�)L\��?�^��y�ϣ��u�[�|e�:>s�x/� ��i�n����5�ؗ�-lh����=����<;Z;*��F0sZ.�1��J�j����<tksڠ_�S)R�j]�ع[59KpA �u��W���u�t��4��C4Ν10��YK�H]���5b����/>�|�M�Z]�q���D��^�ʄo ?�ɠ�o������e�&*��Ou�=��*8��-a�����
�	9�ɜ�DqW�(��ŁQ��vi���Es��mT5�� e�~�%Wm��L�0�h��~g���ȏ�L�^�C�P]��L��R���?O�6:^Hvb����g�ugt�g��{���os.`���ֹ�*M��n }��"p�������\�	���0�F�F���Z�P3��Hy���C��f� -۹�t�iu�_0�����D�@_��e��fˈ��K*�������g����殑E���#���)�����@�{ʕQw�G������T:x[!��Pl����z�g���"�\
睓Xǧ��S�ƣS0�P�`��8w�'�فU��W�s����	������{_�k�!Y6�
 ��S�/0r�+e�<�R�E�e��겺�S�b��G�o3�V�sE� ~c��g*P8A�E��i̍������xs��TA�\���N�HE+�	گ�.�������$��{�iuq�3��8N�w�$�&B��!�(e������i�a1�K�VYw�b�:���eZ�VIv\w�Q�?��A�1igl�o16�)�i͆^g���ՂTq�y>�Tj ���/b`{��%]U����,�,�J�%�l�?5��3� �[��0�p��{n�S�vi���u��n��g���4��x\����q�.�'�}��/���4fHzT`�*��nk������7�g��N�ǻÙ]��x�	�,� B�6��K �,��� �Њ ����*~"��M:��َ���00o�1R��i��>��R
�~݊K=o��0��0�I��j������Lp[UG+m�m�������z����w��&n��>!eF >I=��K�EK4a=���}چ�~L�Z�q��sp��[���.I�Xs�/�FLB�V_i���9c��k�$R
*�L��uZ:��>\��㓼<x�y�A{Tc��K���j���V(��(���G�R���7s��[]r���4h��:�v�u��d[���0��b�ϟDX>\u=�;��+�:�m��y�4�����(��*TM�4]8}`,r�+������u �x�7H�qt����kw?ѱ��.�S� 	��M�B�(P'�me)�꘶��m�8�n�����i��0�����4	}�*��8=n͇�"0DN4oi]WKq�
���S�	��%���#���<T�P[����FS���������Lݔ�ya�R���4R��~ƍ���X}��
�9`j����(~���1q
�t��:��MS�v������ĵga8�S��Ţ܌����Q�v��EZu=F�q�{ZA
+@�wZIr@:��i� y���ǡ���}О�=R��\Bo2��ISzK�L;	���
y���rmԈ�H���O��	���9�ȞcS��6��L�����Pz�cg�L2���46�[��R���O��pr&&�(�XO����)��|U�Y0�p�k�����ަ�Y�� ,vG:iZ����E1n��Z����r�ޚ�l��Kw/�AÏodUXc����'��3���6:��mBmA�r�ш�0�sp��ԣ�nލ=�Ơ>��$�S��7�xp7R$�?+
���<�xz
�XB:4�`^����PԚ���[�C�Q�X����&#���TF�d*ZE�3�[*�����h�A���i|�1��y��e���9��m�TBg�)v��B걋s��Y7��tHQ�XO�wvb��ʨ�|�}f��|�`�,2 ��k�73�����OG3@\�2��˩x�+��W�ݱ�h2\�������\�gc�c]�^(|���������$ìQ�xlH|~X~��b����4�h�g�ݹ�o[�4's!��D=�"d	#럥Ò\�ڞ`�Fڮ�:I)j�����zkLh�I�,���[���S�{�/l�a���)��"�����E�hE�|RL�>���F	 �|�!q��g��'�F@"X���Kπ?�$��QYܪ�Z7nN�v`kO���;�_��"��Q�)`�pC�~}`��=x�ʍG��v;[%���10�,����(K�
ٚ��k�:��d�lw㑰Ϸ���J~3z}��L�ZH�|��8�Cz?�es��۳�a�P*� Ѽ����y������C�,f��
@����"
�Y�w����8j�\n���Mv�b ���^*gQ��0�m���{*���zpw?�ƺ����Ġ��Z��*�����M�`�kf�J��ff����@ռ��_�A�"
ix�D���~����Y��ɕQ�U��y*�m���F���	��MV�r8�+�HQ���{�f���j�?���M����"�j\d΄�V�}���7���S�ͼ�.;w;�! -W|� �;��hb>1�wW���PP�������.��W��3ߟ���������H7|qܹp0���G�xq�-'�6b�C�#�m��=(��<֊�� �aO�D^͉��Ot�W ͆��س�(J	�R�ݔ�o�qo[1������5)>��39��ә��e��J����'��K�x�u���-�X����W��KGv˯���)���_�D���~_��o�T m�`A���*��s��Wa�F'��̠��n��*���7G�I��f�gLřL�������:̵c��Y2���}�L-�q�A�^�g��C�.��ql�j�_���v�e8<���C*q��<�;���g���}�P�-R��Yƛ�wO#���Z�2�½|����s���:s��Jx?������K4PfV��f�  T3�6��عcs�Y�Eǐc���Q�����U^Cjg]ݞ(�<}�+ 7݃�>��"?�;�[G����.�5�kR[��m&�~�2����(�J�� ��嫑ySR��}|w�5���!�K�}Ծ\
M-������Ҷم���w౧^��t��|�-�`��F�GRmï=�h�O!0]��@��m��<?g��܀�)���e1�U�]�A��,J����0s�K���;k[�+�w�2r���z?)����5��r�G�tr<J*U�E��)��<��ȥfJ9Nض��m��b�6��|�±[���aOq�6¡����]�k�d8���4��(&YM��v�$%@9���ziM)����8j�7��}O���]��ԅ����]�U�H~����&���oO:�h��jK_$[ܮN�,9N�kթ������QG '� �7�hj���f��̣��;4��Ϣq�ڵ�22��> 
�D��A~�II�L*�i�i5A��C��,��ߎÕ	LQKf�](ҢF�"�!��Y[� �Y��[��?>̘�f��&���I�$R6�,#軀47/�W�k��X'���Cڇ��O�n�O����H�_�=9E��9���!�+6Y��VC�񸺬혨ʗt0�Y�I���{$ASg�m���d�i(yS�ᵽ��O'�����9Lpl9X���4_�h�R����6i���2ت<���᭎�[�[l�NKq����奐AJ�t8_��#{=��fϐ��d\���tG�V.��Ny��Q.��``��I��w�de�(��Fg��bJi[4��{�i�z����q���c��g۸MW���1t�Qn��6��U"$C�X!�G�܏�5Mk"��l���xm��f1v������z��G�ֹx��V�4��D���s�!>Rjo���V���F�4�������Z �#.Xk�n)���`���m�����/�
g(kq��~H�|�~��0|^��w�H{�
��L�#H̸@dq�>�MQ�bJj�a�S/r��s�k���La��5�����{�e��t橥$�:���\wR����q�*��x~�xoϜL�iz��-���k�[��u�Gb^�R�������T����βm]�I���/�'pW�v�b��MQ���
f�pϿ?kk�B^Z��]����`P�g�/��I��y@����f�.H��=D�<J��eׇ���%4����2 �C�c08�{ڝ�.*��ޣ�IqM��z�c8����ڥ�o�a�>�	ivw��HY�1'�@�����
5Lb^4�4�.�/U��� %�zGR��u�~|ˁN�