XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��*9'�^)(�=2ڷK7XǨ���'W�EN���nդMQŞ�i�_��)���q����k'�/y������n����EfpU�($�B�a�/$I6$�QM�x�n�J�XŃ�4�	�R�>�p�yǎ�m�m UY�
�O^��8���|�O�s>b?��߼Z��C�0OF>��M�s;Ʒ�~�P�s�Et���2���t���B	~�2f6�&MW�)�T�p8�T%��xa�!G�������LփE:J7#ַ���.�w���OسD"v�_<F��fZ�����^�\��6$�&l2�ȶ6�?� P�|��٘�f:�(�qX����46N�t��
S���X�OJ#;f�t����/ؖt�{>��C�hܞ1�� ������N�?G�1�{{6�Q��Qz���	!�-.F�|74Y��ڶo�R���6ل,�M�����!�>f�K?I��!�8Y�%粙!�!nQ�uN��d�\gЕ���~�S�=�?[��i�����k����4�eJ��%>�]]����U��V=jŪb���Vx��[�j/ҹ�J]�nT��|j��-��T��O/e�g��� O[������0)X��$���vPt�Ŋo�m�Y��Q��2P1A�R%%��\1�`2�H����M��p��\��e@�gs/�}��yi��Ƞ��h��r��^$J�h��֩.��z'C�2��?�{�\�I!A�0��G�eT���^$�uy�1r�� 07���XlxVHYEB    1853     810چ��NIT%Ȕn�i�H�a��t�-{e�'`z_��:�Q����X=��>j:� 	/sW|�v8���X�Diu��!'����H��jB�N�b3�W��d�a߸��,�f<��Êt��.4��M���wȾ�{�a?|N�4�y�Q�E�*�c�쫩��a)q��;�M�`c�]��V�?��C4�9u\���9� w~��b��n�Z���c +�x���E�����Zc��B�T��Y��w�i�8�t4��pW������גO8�'�h%wY�9�+������v_Nh�0Ϧ�x�5Sfp����;�kH ��7&')h�[�����Q�E�|�?Fj?151f�]H�?�o�� 3-կ�s���jJ��?����Q{\Cr�n�xc�z�b�l���f&\��@rV7^�A�("BarI���@+y�sHY��u�Ě�n>�<[�g;��]�a�b�`�h.������TȽ�xЧX��C�ܺ �P{q�w�l)d�q�g��	�����^N'	J�����%5C��5>����.;����_��B|�/��?�xt�C>d'��>��RW�B�и��^��Y	�B5���Ğ�,��1��/Ґ��=��,/�Ӻ�m8'��T��o�6�k��c5Q���ݤ�"�Cp\"I9��)�
#�pj���/�P��5K�` k&VK���ҶUӱw����+�ݶ��x4�T4��O���M�s��i�g�p;�����!��m�ȥw��u��e�DOq�� swd�s�_,|�+�	9���u�kA��<g�ځr=�X�"/�����gdTw  U��f9[�X,������`�P�Zv�C�;u��-䚤>���T{&hׇ��wu37Pп%��/۷,(xVbЁ:�70�2���=#�T����FY2kx�  	��"J���N�ً��,ѥ�gV��>��@�� ��?9$�β?�r�˩��%�C�Xh���ۺ�1��o�v8�g�t���笲X� �3IJ�Eh&�3�����ʀ�2��h�F���c����f(~񼅼�g~��� `&��<�hA�p�W��%�M�%sd�^��zP
�)������X������\Ԗ��dI[H��B�*#�Z�?��,n�T��c��[D����M�}�n��]2�w�+�c6�{O��}
n�^nR�=���L=XݴX�g �h|H����hb�m�@���X	w]�5߉i�ܦ�8�� iF�hC�塎
8H	�#M�F����pZ��j�)����3s,N�9��(�;]S�@g8�+���؁B���nT���ld̟���$/2����(;���k�Y_r>�8X���0{�*����9)B}1]����6���9?�}Ϝ�	X'��!.}���Z7�w�P���I�M\��]Ac�LT$^gi 
�B�Y����C�1Kv/"Y�r����=�s
���5j�������1wJ��9�|�d�dɬL�A��xi���3� ��x��w�l:H�U;���Z(%�U�y�uH0S�����>�L�������e��B�9��Ze �5v>1�pA6��W)A�h�q�=��"���f�z��|�"E�oye)U�ұ��B�8�g����)nI�4a�fl�x���B�b"���[��a+���Y�������v��e���" �p�H��͒e�{wJ�?f��F�=�`�����,S�U�]䊚V�wZMl��!%�\� ��#P-�'�|T*Md����*=�NQ(g�tbn��L��,����U��,Nj���U��Ur';�6鋋əuP��u&mF&M�0��i9uT����Ţ�D���q���/�/�!�}Z��R��xaڢ���	��9���E	m���a�T=��B�J�+=�*/7 �����lB!ͮehz��?��������������p�Tǹ�R��.��Bqd����/X�rF���,%�H(�Wi�����3�4:�R\�p)���CD}0��cs������7��T�?9ݺzԊH�ijs>ͪeg��>��so�L�����