XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ٱ�&L�Y��IOȪ�k�9��^o0��^8]":�zw> >VoZBE�_�l��qp��1eS�yO����q��v�ބ�����|� J��!��#��������"uKY��4Iۻ���am�@^��5c�^V��Pz���a�#o�6.�1�U΁�M������6������"��H>�En�?_�^ز�����夎�CX��=i��eX�r�&�S%�e- ������?"�㬴a�G⠲m������Pp�E^I&�l-<�4G�hѶ�K�T�'�#�;V=F�����k�C'3���$��_��5�y��{�R?
U\��}��V�� �i)��+`*�)��uuD�n�=��'&��@���R�:��xe=�W�&�q���XR���:j4�zc�H��p��e^�4a#L9�	p�~��,K@ER����`Y/��R�h�u�f#t�Ȧ��d��� +�U�Vx9�6*�|m��n�(�f��k��>��&�W^��K���Q)����}2�
<4dM�0��8��x��[F��F[$�A\V�"�@'�P�U&g�d2}�&�x�'W$Ht�\��#�|�-�Ѯ�\/ ���� 96������Z��,\soi�D�3�C6:f�����> �\Ưt����}-�-���F������SP:aKT{u+�zq'���J�2�F�@��'��i�2DC��������gֽ��d��f���<�}
c����.oxz�m�jYC���%�Q�j���w�XlxVHYEB    fa00    2040T�:��P�9��C;���O<V����]���p�v��������`,j,����l��)Y9���줭���m?Dfd�ׇ��h��}��v��9<g�9�NA�?`^���M¸��9l=j����0���R�C�L7ѫ�O�,���V�8�W}����%El�h��y2K����v���_p`c"�[%��H��,��y̆N��fjU2
�s�M,�WPf��騀�e4�=��|%M���[� ��v�?,���>۸�2����ֿ�<e����Z�6����=�E�iV��Po��m�G�CGG3{-��UAt60��/�^alli����_�"L#�Z�VlsJxa99�rcp����^ f�G�k*����T
�4�M��&���A�3jѮm�Ū�	��0�I;������"�tzJ�"Z$�jvА�cD�H;�"%3�Ϸr�-��sX�ۿ��xx�o�t^�e�
~*�+��Π���~6��L����CdPx;��7�l�-cEQ�m�;\gÁ��X�U1:|�Z�E�0�	�s�gF�pZ���4�7�Ia���.�K�3�VS�z��� ~p�(�^�c�%A��9R �z�po
��\�1D1FJu��3�x�rL�+1����4$sLʴ_o̴R���x9�'@�U���z�/肎���֕8�2��[\N�ߘ���'�:��+�[.����-��r���hV�\���_�����Wҹ�D���TDz3������!�
�](2��	0��&A%6�!r��b/�]D"���k�1^��a�+*��{�q�J��������Ҹ�kL��7��>!~����fx��M�n$��u'S>(�Ҋ~��\�w+	��k8��W�� 7GC��m�����u,���eeD\��}�_[˨��޹�t��а\Ĩɠ���� >S{�i��'${c���r`⸒���Y�<n�~.�Ґ[+�s>�,b,�4,�oxG���(�_,��i���!��L� ��E�\��o�u~���T�.��ٶF�F�U������(��l��Sk�Y��g���Ϻ�"������+�� �==�u����#�<I�҉ېS����Ⓜ!��	x�����E2͌���u=r{�eҋK8�d}T/pV]O�>kB�$�W�����7sLy�?i����)�iA����1�&p�*&�Л�_��R����`���K ���U@�7/���k��nv�@&E�H\h�Z&\3�-�f�� �b4H5	e��ǈ��r�/�/A��Q0�	*�wz��ʃ��q
�<)�g�-n�r܆��oq�Q�rJ�Yj����
�q����ط��8���޹����'s�Y2F�$䜶3F��eX�6�}�8NUA�3�͚��M��S'���}�̣&����5}��q��`!�x"��B+Ʉe�E�/��`���nt�3	
޳��Փ�įU�zMn<ߙ�O0	2�҈&A-������B%�DW�ȡ��.��g�Ǐ���2p��e��y��!��{Q�2�ϰ7r���O��������2�
?�O3<|�[�����(-9��Z��2����:3�?��jb����߭��5��>Д�#�� �|��~�cF�5X�-21E���3'��ckM�W��c�:�w٢�5y&�t��iVHM�IYs��,�r_]��65�t~�7�w
!+�1�,���\;p�P0N	N!ɕ`�jBBr��r9�*��\�n%�D��=�rŶk���o��a�nS��׏o󻆣�I4���X��
T�l�
s7h�d��P�����{�����M��4�M-*N2�k_b���U��r��Gk��u
�<��=({^�}����Q�lb:�<�����5�b'��+�����a��k�n`��t ����r��QR��`,Xʽ'\0�J�g4;��-��s�[_�۳��A�(�0@�d������z`����:F(�⢥��w&=s�F�/?e�\�EF�[+�:5s�@m�/>FŬi$-��u�97F�+��t���6�i�?'7�i�Y�I����z9%��H���tC�W�4\��./��X:�$�Dh��ށ�ߍ�Ⱥ�/�Xs�Э9&~;�z�0מ���V\s�L��Tω2�dw���b��L���u�s�ŉ�6<�ުmbu�)]��+���"��L�D��.���������t�p���P����U���W�	|o�L=�����N�UL5��-�*G㣤�C�l�;o���Y�E�a�g�X#`�������#�Du�q:%F��+�2�ɶsE�Y$q�|��X2s1��P���i�qRE9'r���z=׏�h�B���0]�6�T7�9An��}?��3~@p���[Jj����5*�O��L��-B
@joaB� ����,�ַ�g+�ɧ���cF1�b�o�c?��S�\I)�Y����_��S�ǐ�6e��љ�H�ʠ����Jx<l�j�����������zQy֌�&�<WL��_��%+PM2��w�\Dƫ�c�S?���䂊���G��O7E吘	�L��R"%�Jv��pQP"��m�����T��6S�gG�1~�pΆ@���IC��kU����2UKk-���"J�՗����� (Y.4�6C/F��Ku$8(��ά�'��^���2����!6�%�]����Ȟ�������% i�'��<60k�|1��/=���Cd{5��`�'j�߬8_��4Ep&4m=����UifE��(A�H`q�[c�5��6�.��݌d%vz�@��AbՇon�x0��vuA6���ή����b��/�dw>��H�߅���_	k���O���y�Z���%�D�n�#P��	�B�� �Tq�ɔ��8�G�$t���M�M�є�R�t'�\�9�G���~��Z���U@�}r	��?����ָ�_aG��Z
TÆ*�����`w�� 5�)�.L��ߒ�Q6����2B�����y5���bI��4���/�CK"����Xi�5�9����<R���s��Vl��f������+�,�.�`z��)B���i� ���E�B����AmR(���@���篛r�ݘd7�j�ka� /^���c��K�����u�(���*�OlL�2���<)�ޟ�R:��G�fk�4��[��,��]̎$�C���t9F��j	��I�8��͖T��)��d�*.�'�
A�� ���w�g�{����cuzH�,�W���fW�X zR��Օ�
%?������F�ɾ4�-�k�C�G"�y*�{���2
92�)'�(�DwZ�~Y���:CQ�����':�1w�@�7��3f��&9������Vl�)׾Ykj�bosh�Z�2���âQ��
�t��MB��M�	ZG���n�����&P����U��(�Mf��_�K/��pU9�!͆_7���1:�_��@:y]��6����p�l|�
�aF�L�����0�h���ն�<;$@�3�
�d��c�*OS%��"�(2~��xE/������X��2����u���|���c�H�wg�{P�8B����>yA1����i��_��(r�oW����w�Q�)�ˑ}�rE�0	G|3���� �!T�"���`�>XPj2Z�Ď�M���L����ng�}�2�.�"�Ig�N�=%y��xVBZL]0L�6�ܤ�����]x�Hd"<`O@	���i�N>�?>�5�ŪF��3�Q��~#��5(���`�H�E�os���D�V|���]w�M̈́����v���4'�ֶ���w����l>�7h��_�	R�b��T��*^$�����DY1�I�dp��]�E�g5cƳ'��vɮ�we��7U���Q�kl~���R�.
 &���F�;x��ӷ������2���Ͱ,"��M�O�q��=�!��sQ!�X���6���3?+�nZ�Dk��'���:Ǟݵ��є�k�/�=Ӣ�T��5H�-R`r�j]�n�)a�1���\�[g҇!ٽ3�"2^�0�=�ȶh~B7�����/�@p�2�����#ѡ�+��eY�d��u~c�%�(߬��K@]�s�t}=�Ā���-rQ#��t�!���3���68�P����w��䜋
��@�����G�I�����������)�W��p1���P3�k��A�g�z�<WcVےX�8	d Y\�`Q_[������w(` u������IWB�X8c��w��.���o�������ح�"s�+��2~�N'��������m����Lj"M��'8eа0�0&�+�t.��X�Ec|�(��O��B�3�������#�њ������<�;c�w2�%>v0d�)ZJ��q�I�),9�b���vhco��]6'O��[j7(#,@̍ר[�'5@C	D=ى�����2c��w|@��^NWr�M���y�4Ή�n{a��7?`�0t�"!u�&9@:�=Z��$�*��C�udΗ��	�?�0m��?K;^�J-�Q|���R��Cc�Ҡ�h>�*(/��`ȉ� W���.��j5��!lH�h ��M��[bS�u�K���������	^Za-�J�}�
��u��צ��$�
DPT�v�p��^ѓAKƣ��BԳ�<��3��,��/�x�����r]��3��rQ�������2ܘ,�okM�%�(����3��u�A���0��{�JK;Y�j��1�Qqg���~�K��֞4�� n��:���0̱%k׹A�B�ȭ`{�^H霽���B���ٰ��DY��L<B�V�$�`A�5ӷ	�¼�7�f���d����4zI�r��CF
~KU�1v�Օ�_>bE������}���o;��*Q�P����6�tY���R�܉ۘ����fx���.��O���_�H�.�PV�E�"���/X�WPL5��=�yi1���#�����5��r_FF;��X����6;p�y`]��C���h�K���-�m�J�ņE��9._�}
�+��-PpPe��n�[�4� y�ǝҟ�2�젫.�>��;Ɯ���d�,g����B`> =n|YO�T����q.j���g��A�������|�/�ewu�B�:|��@�n�c����G�q�Δ�_��?.{{�,�pv�'5���R��� %���#�rz��
[l��|�����U�d�n$ %�O��2V���N\�����~��^�5�cnQ����A7AY��$g��7jte��Q�B
)B���x~j�bL���5���0 �QM�s���B����yu��� 4gA��6�E�g���i-zG�pDo��#�i�Ö����#3���Lk�����y���
�7?TFI<_6Ǟn��D�9QXG���wPt��c,�l!��!�K eQF�L{�bQ^�yO��Z��}��)�"�ͤ��\T4J�&ˡ����G+�0#κ���.���J��lԈ����9*�L@4Ό�f �7ڽ�����[�]��tě.U�H����8��ƒ�Fr4��EE_݇.m�k
���
t�:N��6�A
�¤�i�9~�p��t����bQ"�Ꞩ��5�.�aG`��N���"�P�	$ GS:+ʳ��ԱO��S�!�H*��Y�.B;R���ߙ����16:�z>|��#*�+�A���R�����^�j�+�^����?i�]�в}�r��p��_�&�MMT	f6���]���qg�"�*_�<�D'�:I]�~����GCE���
l���q{J���|ٕh��4L.����IS;75'��B�%����S��Qw �4@���t���i��+p2p�FǯUT���	�-�li�*�!=�Nʏ�D��3��tk=�Y�y&���z��*|��ƅ��`���%���؉08�rHi#�N��1��f��K��Ӽ� Q��:�����!��?ri��r��͸[��-�`�ԜF-2e�m�k�WC>����!����c����F���y{�0��ފ���Xީ�a�>�8 �6��ֳ�4�%��G(D
�/�R�㖺^�����7�tE=w������:�3�|�)��d���{�4b�߃�%K��{��д�.�/V�;[`�6�>�,�Aʅ�yR�����ri�Z�+�� 0�1�E'j��us!��Sc��S����p��!�q[���S���M���H��-R�Z�uT$2t����V� f�l�<;:H��v�/�Q�W\�CK��F�k��[a�A��?���>���fΧ�Jt �@�
m{۳�z��;�㟷��� Q���s� �(<H��m���������!�P�8�q�S���q����kaAmDD?���K�'�#�>,'�$��DJ�4#k��hCdwen�2Ί�y-����ݞ�OxES�G�;}�^���w�Ym�7=�=e]��{�'$p��=���1ogY�ۧ��MFb�-�-1N�13v��(��������	n:�c�珷@�J��k���Q�cS�Ut�b&�e�V����8B�2���bH��2��� �����"��G�x�U=�Rs���٣�?��2� �E� m6��Z9|n�岡��h�dP1DЅ\^օ;��7�\����,�q��/,Y�}1�ಒnfDI�OE����� �����3����`t�����3���|�T��j���a������9݂�{$����G�0,ؗ�,vC���p����L���!�fD��\יQ3�	�{�9�G���e�Us~c��8D�=W5˿�L:K��F0а�o�	�7d�ۭ?Msl�P�zۡ\���F3��(ey�����Ȁ���r�Lg>Ⱥ��p����U"�\�k�hi���S�A�5�b��bCMd ��:�'(��HV��2�]W�Ӷ����[ҧ��g����p���p@ۇ�F�N���չ�y;�%�|�&�Oy���S��POnBN�VUB����$P�,5�4�!��J���3Xw3��L��n�������OZ��Zƞ쳼j���Z�%��!��4R�f�������'��7���R�?#缁jI�G۴�7�e>�֒����)'����� -���z����e $�����Sd��ؑ�LrHC&�����p���<.� ޼����e=%m�lL�xj�o͚I�D��&�$�ˋ��u_��͌��0��|u�R�һ[�c:]pAB����>���"uPV7��n��uHo�����!Ap~��q�8���<0��4zgH��L
��&�҈M'B�*R�7�>����F:�4��5��QhК�~徚|V��f��b\ƙ��@��A�$$��y��cP�h�P�^d^k��G1X^�j�d�dM��<�b!���z�/"G�i��P落�B��%l^�x��G�NJG�-Q�j��#|@|]�3��ks��d3��^�� 1`�S�#��i�hE����'˦;,�Z��Z�z,+�-�Y�tu�RjV<0�p+���Y��_���ݎw�q�C���_�J~Կ��F�ĵf�E/�Y�L=���ٲ]�f�n0��|�!���(���z�����Y��H073���)� �
�Q�	�u�-4"8o�d�V�78�;n���3�{�AH�ek������x��"8����5������Rv�kk���T	� �y�:������Wnpdē����}�6M�E��y�R;�i��X��S�+v;�8	f�.|���͇��)���Y��W��y��!���PŤ���4�wR�?Hޒ���I�\`֏�k`�뇻QS�#D��0)��#7��%��®��2�`��|�j�N���N)��^w(����Lҧ�ˈ�其��ܼ�--5JW��a*�=��u��d�qQךR��� H��m��]:��uRۡ/7Q�gL�R���4ڳ��B��&5<�������gl�����!��2�q�Һ��WF��>���¤`�f�R�Z.5?O���g����|������Iun��x�s�ļ���q�N�<-�s<k��ZԼ�3]��w`G&i>���K����Ĕc�@ӹ��L��:S,T�@-�C�OVMJ�d�8u���	�"wYd	̤�Yk����B�K9�|�H�XlxVHYEB    4f62     b50���7�Ja�����*�C��퇲�*~5�����]�c9e{�4�Xӊ�i�H��l��A�/;Vdv#�/]�^#��[�ѥe�j�w�U����M��RƎ�w�.6j~�����h�����
�u����'������������ Ƽ��R+ӌ��#k�"��'X���"N�'�����4LJz
��h�Vp�����I1	z��/V����l�M4��oxd��6�C��'�dO�d�Ȕ��TU�,<8Ӡ�hL�s��;pO]��j���[��&ϞT�$V�/!y:lF��iީ$ޖq}��F�X<��g�k�����'�9Ls;�A��7�[����ۘ�lz�R�Ӂ�:�B��q��@�X0!���f����\��f/�&!ߘ�d:>/�|R��^���3�gj�P_�2�(j�B�ҟ��.(���NDܑg��Mi���ð� Y��S?nE��>�LEІ�ؔ�-Oy��<�(�Y*VnZ �g��{D�BQ�QĦD8����u�Ge��c�ӭ������)M�i.]�+����,_�ҖY(He'F-�b2�biLb���	;����+aô�$�C�P���R~6���� � '�AGn�]�~�-��TTNӗn_�S<��:���������H��2�a/R���i`9i��m�[c&����߯�Zw� �3&@�]-i:^�'x��M!�D̬�����9Ã~��[��Qs��[�¦3$�}M+��nr�-�;IT�IE�Hs �YҞLZ}��cf�ۄFh琄I�S�u>.��c���B��E~��2~�zؠH�)�e��~��YYA���޿9�|��xl3�1$��\�t��<-	.���,9)�k��兌޸��u� W�����'�䡮%$����D=��jU�:�ݬ��Ag�M�,��*�k�Yg�G�o�L����+���ڐ$O�뀁p _��I�4�W&�zO*<,=�:Se�1^y��:֬A����-�n�_4h%�U�� �"�?U{ �Hv�����\�	�uT4,u?�Y�r�<k�5r�j���̈́,U��M�:YA��Cq,��P�
ً�gC;�f��GGV�R
ln����4V:.pr�\��?��K�j5�ަ;�&���|�#�>�=�`lD�@
yv�C�6]9���X��U�Q/KX��us44|d�*���n���%E/���цru2��0�F�Sǚ�T�=��2�K�����+2�9E��^�� a�����U��&��Kؾ�,�q)G�� ���&�Ea0�BĪ�~���B��5N�Ww,�xt�:����[��I���bE��Դ� @��Gc6�[.��{�HvȎ�����190e=��]/�w��+D\�c�����s,�����2~���ؖ9
#1����;$B+������d�&Ӡ���L�Z���o�O� ��3Z@o�)Bh7�<��f)"�h����xF���1��߷9��;��ʋ�����?�+�n��L�;=
�8���U�Ďe|�C�O5�a�R���q�ޟ^~���)���yB?�q��s2-��7G�gޭMH�Q���$�5�rHʬ%׉A�(��̻�����IW�R�
m�\+}�bIYzjԍA�d� ��V��������̀��픃�_���b��4��M;3� _	��6!�G��+���eת3�O ��,\�1J�/O�,E�e�!,e��(��#c�1�.�$_yƼ8�Q����E}�R%{�<�(P0Q-�m�G�n����؃���~�)�s8�BB�Jm�2#�Η�g�u>Ux�5}�C)�~������HH��j۾����j0������T$$||]��\xޯ㻄{{�����::P��	?�:��[��T$h�����2�$�r�-c����SO
<zQD�5ߖw��ٻAh�`#���p7˼2�Ї$�5d)Nm�~̪� �>E�'#3 vDf����qO.T0�o���7�O'�&3�H�$��X\����Fmjj+�HZ�fM�r�u��g�LJ��G�>����w���߼͟$�غbD��b��=�S��V�3�n�:��8�r��I��ֹ�zwU�`����R�o��T�lS����u�A �;��`�Ĉ��Y��h�P�׻��t^��KvC�	�-���3QE�a�E��'��ڡ~-��]c��bٕ�dƇ}��P���"ti��� ��ߚVA�Eh�hL�1�~=S��X�JHM���E��C�����E�ڸj<�r�9Ҁ�t�F�P���J�{\��
�JoH,�����Q�����P�eșO+��b�y��TJ��HEky���Z4� �%��B����W�r��z���rҋ~���Щ
t���DL�Pp����J��"��8s�	vI�Gm���֩��M����ՠ�[HƗ*X�(ˤh��	��<<��"Zc=�h��V����L��K/�)?���BKB��"/1͖����d e捿t!2�P#�E�r�|����d�+���*$��š�aWy/�e��GR��ũQ;$U%�J�3�����P^��5K��Q%�ͭ���F�8e`w*��@�ȧo�6�O�Ũ^���e@��N�:��<%�L0p�o;/�L�ә�<HZ�)YXܸ�8�+����&lO�;b�c~ץ�vc��s��t��s�0]�A������N٦W��w�a2T< 5
q¥C���޷{��?u��Ŧ� ���X�Ԅ�q$k��L CG`�'���Y���߰腏 ۥh�Z�֖��M��)��Rz�������P��ф���~�Y�0�/qg#�.�V��U�1?"���kw��*��@+�j��KyѼ���(�P�]��H~�@�tݎ����,Y!/��Xќ�8�z�\v�8ӿ�^�