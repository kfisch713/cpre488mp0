XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k�)٥D�x/��5;��'�ZM���McZq��Ӂ�U�Act}DT����ᬖ9Ё|�,H�63q��F�*�Oy�@���� z�-����$ ���Бza���~�l?��i�F�uQG���{�<��+���Hΐ�1W@V?{}�w�|P[_�wq�ϣ�P���c�|������% �7�,�E��X.`�s�N`�!l���Ib�Ff��$��O�ef ���9#�;e���ffC#���;�����y�}���Zzx�7�N��)fFnN��	Ǐ6)������dC>��¡������۱�<95E��JѸ�P�;ڕ� ;�
�t��&��;2ÅF��E����趯��AJ�N��T�l��}k�@�5���7��kO�xƶ^I����,�ź�����eO8��(P���g��s�[���3�N���5�JP�"1'ּ���ٲq�i�=yXƣ�֞���Ex��Z��uL�N� u"�����nQ��{�5��*X��BL�!��:7[�����R�j��z'���<XP�gEΖ/�D\�ؖl/��.U�yG�<�`��ɠ-=�~��cz�%Lj��:�WcH�Ox�����>�%.(���;s�����4���h��}����?�!9�D�Ev9�M�K��b��W��Ii��s+��`�4bo{JA9�h��O�r>���_����|��)l2��!7v��H�*�K��Z�Y�A�����w0Z�?�0p�3w#P�R�가��;�v��¼Q*���]h��v-���)���*$XlxVHYEB    6014    1840㍀#m\"r7�$�\�p��]|�:5�1m�;\�a7��|	��;[K���������0 �޽Y��$8N��G��Z�
|bq� s�Kf�3���o�A[�]�0��7�*Hr�(7/���pJ�rU\ˈ{X�����]<�E��rmN(Į��4�]�<i{�G����;e����8et;�FY�z��pq�+6TIRoK���c�e4�<}W8�"��)5	��_�f�u.�#�- !a�E�Յ�����	V�RF�(�������(�����$猛�y���@r��n]"ņ��vr[c'V��̓Et�Iy��1w>�y�3�$�'�f���I~-���Ff�sS�]ءU��"��2ˑ���#0K��i��W׉e��j33�m��)� 7R�*@o�c�"R��&yRG v�|��.�]���_�TfU�A���<�!���k��c�{15Bx�ن�#Qx#�ݻ�
 ��U�v6W�%t)��$�4i�H��jU7����Q����$��{���_�c�v���g��h ��m���[�W�4i\l9%z�F=H�2������	��ۍ��>��M0���o�.#��>�f���"��z��돫R@i����c�8NY�9}�����/���1=�������]�j�;$M�9��O2�eb���7/��hΛEpnUJ�a���%�+�$�J��s[1�'�O�I�W<!��@���0DM0e������3�#���?b
�"k�B��jas��׌ʼ�P\��ʹ.��CY���2dNg�Ɵ�9:�zB�;c+��o"Xn	�Vk�w�����$q`�̑77��>8�&ȕ������o�M� £����}?Z�@���4�� �{�ך����>�X���9��˗��ڋ[P�n
7G�6��Ũ�_��:���CN=@Ї�]�q�Dw:*�(wt�\� �k$x~]�R}&��5I�5;<�4^�&��uǍ��C����:\�KI�X�*/���������wdB�Q������8��+�d����[R�{������[�l���''���}ȓ4;c��c{v�T=\Q�}I
϶.'��!-7��Y�g�O�,E��h��ޜ8k�ր��>�(�����h������)��շ _~�������|�H�L���>�x:�������]�<~<wm�\xJI�lg=N�f#�3�+hMW�A
�SY���0�d!���_p�=��v7K[�n�FN��:��l�R��)K�v��$�|�Դ�� �����g��C� �ʊ�L����o+Lwkf�+���9B�-e�E9׮�0�V@n�	��xt���V�gN�nPǢ�]#B�ϊ�̗����M�j>���{�d��-GN��d�NǑ��M	Zt@�5�ŗ�ئ딦Z\���oɗz�/�N�7�v�+�ImOC�[��Q���V�ԯ���T�8���ō]|� s�B��SQ�oۙ-=�Ʋke�4�9�e��_�LdgfKx���x�e���['���ӟ�ߘ�@b(��Sԓ�]�aI���ux۱�����G,斦C׺�Ql%�������`�l������i����9��$�a�';��c裯�u>MҧWW0E�$�[��������l�/�p��ݐ��B��DS�h�KA��]/:�X$
/ID�7v�:�u�K���ʥ�)�=aP<U�US�w��<2���=Y���N��<{h#D��a�]�½a��-�BK�����>Ո~�f�y�T �/i�El�� ��/}�KD�q�Wp,^�"{��e�]H�l:l@v1|��A��XXz<�4����Kv��1��I'�Հ��,�}���(��c�a�����z��#�#�8D�񋝁�WBB*'i��ry�0�(�;~e
$b�T%��e^�"���m�c�s#���u<�Q
�E�����r`7Ⱦ��*��n�����|RD`�w���L¾��]���d��eN!ut�h]�6��H�0ߚz�(%�j(>S���m{��8U7v�-u��s�` ��&{��ꉚa}_\�x&�7*a6��f����!:����a�j��es����n0�!����N�U�LC}��ʮ��JRw�?�JU	��O	�u��^da;����I�$_����oكaCCd�̗�(Kj���j��Q��/>�2{O�����oҐ������oy��&�E��#-�R��]�/�ũ�$ДL��a3p�ݖ�������]��ȧʷ�9����W�}޻�)IEς���f�A�V�: ��-���9�ߒa\¢ڹ��\~<!a�q^�X{��J�p5I�p�tl�����9e7�b�NfU�-�&�������(��GJ�q-nQt�^m�g��c���"n̋�3Ah�_ܠ+���� ~NӴH
GWׄ��`<e#�qU_�U:��l�?҈R�U/u���MS5�r��W����JW����'�m�i�\n�^fU��t�z��z�LJ�L�u/1%�n��৊o0J��J�M�įW]`Ib�c&!Kq7�`�3��}�Fo��DV�ٛh���SHjW9�;EE�'H���/E��/�~>'�t�<�t�U���Pd�Q�����k��I�"b��ݑ٫��7�ፓ��c����U�6�9�'
��&/X�����u\35���_�}�:bX6��m�C]P��0s;G���'ۗ���MU?���^�pu}���\�6��H	 L{��g7�����	�AZ	%D;z��;�k�.��Ƭ�F�����/�NL�@�N1�BC>@�A���[��z���v���Uk�����J��9��u�G����f�z��	���@{�X����X���4���F�p�3.�I����'B�5�"�x�U ���i�r����w�_z�M�f�̒�S;s4f18��F�'��̀��S^{�fƿ��k��t�&&���L�#pN�3�4	v'���X�Ob#�d�.8X��ܑI7�I5�U5�����+w'S%������ta2�?%hB}&�i���:aa�Qy��������h>�z�',�����^
�������H��`�D�J���Fu�\	�=.<��=������P7E����~�x��s�4�O�x�J;Ưn5�J�����-<���[ϛO��=6�����.}�6�)�0�7V@�ְE+Cɥ4�H�iCo��I�g�`���1�5ܠ�F|� "�",+G�-N�����-�o}33�Ĳ�"�ɏ�6��<�H'�*�7uK�Hc�+�?p��.���4Z�N��[t�����8�"��%PQ4*�>1��y�g���9��y�7�7j��̓�����\�ƽaN�!�]�O5/��ݬ���f��z�[mj{�%_�~���<$X)	�����6��n>����8���+?N�7�!�fQ��c���N@<����E"%����=$��˟2hU��K�D[�鵒Y�h0W�H|��f�+�z1�u^�z�D
cR�k�@!���D�c�N�]�:;��:�9�D6��\$��p*�X�6X�z�n�V�B�=CI=�BY4XpP�,�͙/$�Gc�����D�IUb����X=�x��DlhɁT7�8-
�P*~]"��d����?�y�y���~�j�Lf�v�-&��pu��sY��fu��(��jo��i0�U�K0J����#Z���dX��l������ۉ� ��y����������9�c픗��Lv�c��q��(®�N��M5
l
�������\���ϸ|�Fc;m[28M�]\��vsg3Z �S�8^��-��w��&�v������r$�+z]7���������z� h]:���aa�S荵�%wO�yKʢ��e�tC�(ג�Ȏ�Ո����Y�x�}����y�`�P��ȧ5P
���)@er�ˢ�2]4ⁿnd��G��L��0�� *9�xz)��|����X9�`�>���TK��L=�:t���*Q���#��J2 ��#hs�iT=v8su	�y<��&t�����B$M�=���mS�ڱ��ar[��( Ɯ��!Zv�<_eK��:-Bs�.ğ��s�a��(1_�����_3�֟��e������UY|Cc.�*�݄�WR���&PM��svO�O���H�s�c��'yg�����y��[B~�5B���Y��3M�QOY4�*���"7Uױ�,B���uT�bHT��=`{Uͧ�{��%:a�j���T ��k~�叵 6�QA���Ŷ�|�`�V�yG�Y'��LEЇ�;5Pp��E�;��~���0��Q=4�.3�(�==���V�	}��R��,���cf�&@A�߻�Wds�My!H���,.��;f������A�}Ly��W�{�����ZB��&;\��3<M%k��ue=QC���g�ԩ|'�t�/9�L�������bkk;[�'ҷ��ƃ��?	��v"� ��e!N�rkmDy`��ޞ!k���!Y\�b4$�a�Mc�}�5��F��zD�t��v[X�����4�%����*�H UfQ3ڻF�iR|��Hjs~������@p("����4����K>�K�}�6�p,QJ5����/��	�G����Y��+�M'.B�]h���	�6#��U������#����H� w��?�z�獯��/(P���H�?1�9g�@D,T%@֌�4��!�w�!���1��X��F6nE����kϽ(A[��<=cQ)�J�y��)��P]��������,3����*��l�E�EWY���P?qB���<�e�@F������2h����Ã7�#r���x�q?��;G�ؿ�p��^A	�����-���E��fǾw6�CkԿ�+IW��B��	Mp��,� ��g�<,V;���C��o�n�|�0Ӿ���B��;kD�+����ۀ}�P��qAB���x���{VB%)Ђ�xHg9�d_���E��n�SW�
�U��z?���gX���
��]>q�����~?�önd�뉮���=4�����7�<��t�X�tg����C�Ą�57�	��2O'QE�hڿ砗s�M�a�qI�J��qZӉ�C>��� ��u;.���,�E�R���B��2&�iʵ%�t��W4_���1�S��zu�v�O�3��8��R��ߠ٘BdC4��z�w9!ݏ\���i�-Q�c�д�� ��W
�����2��}��/P���xpӯ@�Iz-��P55gd�7ѧ���]��9L��Y�ȶe�u��W�u�I�������
>.�Q�ryb�,������:��+&������	��'{n	��ɤ�5�[����c�W�����g�v����-0���L����֗�Ҽ$%B�ɣ5@�f�f�$�D���|��	`݇�SWc��'�gb"|nz=Џm��IA$T�"+�jb��V���5)��d�5F5��wN~�������	?��S��D���Oy���YH�4�s`�
!)pN�O�h�ZE����#�aܝr*����?�3��m�X�S�����x#Z�JU�����ˇ���kyA���ł*k�i̦���ֈ��|ӛ(� �Lx
CQ���$_�.� g����M�+ ����H�;�I�Lƥ��a��}:pGⲫ���:���d�`�5��K|�2�C�Ф�7��f�t�ud7��O)�g��� O#�P��`o�QX�Ä6P�LѸ����'S�+%���Ӻ�t%X� ����Z>�NY��(���_&�έ��e^��$؍��qX����28�:���l�r;�@�����ԏ�؊�.��x�[�6�p`��Ct[�E��5k�JT�fkg	�R��	.X�b���ԭSoS;��nT>Pa�JT�m�)��Wo_�]�z;�7����c��AHQ_�%��d`�[c1ZV�c�Fԅ��G�d�"�o����Y)TEAc� 5�Y�
���*�c�U��Cޞ�`Hj|��r,��pT"�\��$��5> s/�x��+#�$���+,(�����(�b�Ox�Ds±�_�!t�{<pm�ц0*������(�9�"@]�zgQn\9M�@�j֝�q2�4���;���MJ��0 �-sgE���gsܤ �