XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���H톿>�<#�+>��8��>�V�O��,WpA�iW�g�k��D���{��G��c���[R���L<�'��~3NŻ�l��NE�oK�j����Ԉu$p�_�<�93�\X���i�ܨ<�H���y�Q���P�y�d^́�3�c�(s����)5j�"�	;�v}���?$#��5r7���X������iIG�т\R�jK��w<��*"`�T����	�l�
S�G�ɾ�L�0b�@��>l��1޵�i
e*���e���.�1�r��$�r%'�H�}�pY��Z����/?�o<��Ri�x�A�P:T5	r��4i�/m�^G���K��I	A�gN��Y�;���h3�.��,��rܜ��@%o���$9$������n�@��Ke����Y<h��9%�����Ny�����s�!,��ܐ�d���r�
�Y��� ��|��cli�L��ǫ�Ҷ̚t��΁�tjσG{A�6�궃�CF���7�Pʷ����
Hz��c��b��&�-F���(q-V��װM�JY����'j�p�a�}�a�հxH���li�����6FnRzX,�=X����H[�!����f�ck���z�v@�[-�Y9��n�����`_i戄<5���y��O���ԭ��F�A�Om����Qd�B���YK3��uP$���[Nf���q�Ly����q@b<խ�O��B�W�՞�:�a\�']���uFR
�2G�k�?R����3���Ն��������� XlxVHYEB    a037    1fe0��̊��M��[�}P�$�Q�]~�eu��BǋZ���bѬ�gGfb�ݙ1&�<����>Ae�)�3�a?��1��E� y\~VO�S]ϖ�I�*�~��6�=����o�`���7��#ƶtj_���SV���;�)ݡsruF��Lޔ�-6-d�$^�7S"�^�t[�rn\� �C+p���
��2ѣ+3����ȧ�(�H�3���~�t�n�� ��Ö�[��w�Z����^<���B�����ӷ���;1o��.��~
�B�u�A��Νi_�/>]�ĦP�I�q��VG���.{��>;�8�J�$��2(��\k���3~F�����r�&6aC��Lb�x��iuE�"�)��£4�jy���\�F�M�6нf،qUl�q87�_|;���++e_��>�3���B���W� ̫*�έ�S�X����$(/������������{s�`҉���x_�P�Λ����N,�����5p]�U[��g�rME�S��hR��_
��Ef��+GC�������n��X��W^w�w�
.A�A`(鋌��NX����8s�y��bB�A?�v�)e�d&�<������й�$%p�"6IR:��;GH<\����Mlcرs�T0�&,�qpV��W}��`��e��-&+ګ���1j�[?S={MVN�S���~�vc�|���:�T#�*������?��E�etY�<n���y{�:�'�c߫�0D0���IYL�z�!ȯ$k/�^=gW�:K��m3�*gjyt�>��d8�r�ݘ>7Uc�a�� ����uf`�)d�%L�C3NA�j�]��CY���:�1e�F��Sh;�M�N`)��W��#c�L",�i��d�jc�u~*������xL�V.pv�O��yKY�3֔~����,�B2/A�Q}7W-�D@�E9�?�E灉"�%�3�	[o�mI�] DVf_bбI��?{3_�s;y�/P�ь�#]j7ouy�����&!�i��n9*�Yf0<���b��[�<�x44�'�D��@J��vauW�͐.�,)j�m9�&]J.*��i���S�������Z���_N���s�c��R6��Ʈ�v��շd���ٰ�Cc��o��e���<O5 S�RH��0j�~�/��x�������(��Ĩ!�J�xa�Z2<��y�G�KU�ܒWL�۳҇�P�1���O��!��1����_t��K^;;W����|R��1υǼ�R�NʯͫVLT�u�[3��CC��@9�H]#�[��h��	�~j��&E��ˇN��W��47>�R�X�Z ������r/Z����A#4�4[g�Ư�h����ekKr߄)�V|ō<E`+B�#n¡�v��O��� �[���<P�TЄ>��9��ǲ��m�A�᧱���ï`�4�_;�MwJ�d{�F�6�6������g���<�/�W��[��($���܏I���5p���#d\:��#Q�3�`,�*l�J@C�{>g̶��5wZ:�h7u�-�F�\x�ikk�%^+:��k��'�Å�3�wVO�s8ObV�Zis�!��y������m`q^FSp��<ϣ�`��*���n�B3����47���i:G�p�O�w�=�l?+���@��
xՂ��Nu�+��?������S�A9-�ں�0$�f��2zR��I��e5U����7صc�ȺV� �C�L�I�YYx�����Hn=�4Ѯ'�͚K[��鴞��Kp>4!7�h؜�Ff��$y0��D� ,�3��i;\��� �񼽶����3��������f�QB� +դ%P�7��gDK텆��
�O��?f�S��E 	������h*@�������v�#|r���HO���<�1���+�oui8�"��$�PX��l���1��E�N�J�W�m���1�=���_ ^����w���9p�9ˤ֓.']��T�&�}�> ;�g�4��s,�i%�<�<c�&,�=v��{�#����}���cH�-TA
�7/C�)p�M�>bʚ|��>BI�t���J~'^!�c7!�L����G5���Q�����i5�&Ď������C�r.�o"ތk`S	3f\_=��8	2^��W���:��W�]I��p�{-Ѓ]�sD��y�*�Vi���+�WW�i�CŠ��%�轅��>�!<�@�H���!^/�ԛg��{�Y^�O��TB����	��Z��<`%oG�Ծ��- _��u�f�d��l�%3}Fæ��r�v`�}�C$@e���4��X[o� ֩����!j��.�\5b�CӤε�E��͠C<�[:m��s�Γذ7h�?��j���RA�L�-��!���N?���~⳯�q�Ee�F"�\�Î�7�%٠��aHpa�{U��b*�s����o0b��$�����:��5�y�w2�=���Q��� ���ߖhΜf�J�3\��&W�~�C�[��V�����Jwǩ�k�@�	��ǎ.��j��c�.���Cﮍ!��_5z�E`�>���������!�M9��gȸ��i����*�(��i�"���UΟDn�%9m��3rj>P�L�"o�MVs�C쩌�r��{���{��_��0;� D:2I]���a�Ut��׋��C�sOE�1���P������-h,��$�$1 n"�FP��|%U�!�G�R��~������v�&����HƼBJ/t^�>)]�':��{c6��ݱ*� \-c�7�zN?ˍ�s�l��rXԟ�!l;l���c��,e��?Om6ƫa�]�TE݄�����8ʋ�Tήmp�v3�㾃>�o9�Pą)�A'ƫ�t`=���K4�Q�\��4�9dE�O�����C��y�)B�<�a�4��qky���N�D��%���D����ǹ�����M���	�A��vW��R�ZR�:qR�|K�f�����x�g������h/�eaIn,��� Ĺ�v�g�t$��J҄w����O�0Դ����\+��̋v(!���B,@��O-���We
�u��H��7σ�}�.��!L�q*�����uƚ\Ƨ\H�#�Ӏ�fNf�҂��"�G�q�e���$຿@R^�}��Aj56xE�p���rn>�6u&��bt��#~��p�x��������~��8jn��/���� �@&��련�J(����ѷ�h�jX϶�7��X�ĪO�*��(��<+x�?1�v$wm��%�Y�L���߷qF`B%(��B~��vB��g�-j*nnFg�i��k���f��p����	]�2m�rn��HE��K��2y��mB�=��*�x5�l�L�Y5���Y(l���A;dn'.��]�Q~�F���E����#d�冩�lp��[�4�?;�	N����l+ן��&�aQ]���<Qm&Kn�ٸ�5�S��T��k�sm����!�R��L=�.�t�D��I�Y�K���%#�V���8*RvM���k[tt~��N�<[��s��(�7`z�=�r��I ׏���07tE��Loo_�4��ً[� �a3(�p�����u��a�T@j�D��x�I�l��'*� ����W�`7��)@f�[RΏ=n�qo��ղ��q`O7&}8�a�t�����8]i$>�I�,���@��o�$H�ke���*�(W�i*����lOy��)t����˛a�Mfd\����O�����{��R������;΄�I<��Ҿ.Lm@X��>��T�D�	7q�^����sk�j.˾s
�	��&;~J�e}9��͇q��A��u�~��6V��7X��̦yZ�W���Y���?���> ��k�i2��8���{*͙8K��aa�����R�:U��|X�G�Wĵ���o%���7����a�%C�AV�4�$���Ս��$$'_��a��˰��Ƅ'<�r'y���~��͑ȹKR��g�v!M0�>l�
�.���{���� �"����W{��GRx�S#V�'G�R-�U��׋�7b�Gɶ5e�F��A���Hn��(tk�nOCh����6�*W�8[�l�u�b� �Fk�����ʚXwU�s�gz�_ɫгߌ��!�t��7�3�g>�L��m�,���΄�|U����.J+�RF�|�v�A0������>� M���z��{y�r���h���Zm�cQ�VV��˳��B6�:�[ �ɐ�)���Z��;�D=8��:���(xN��Ǽ� $�5 ����_��A$�/7u�%����Lă�T��|�� �NCPXop��5�0�������_�� ^�Ǿyf��.���4,�(�g{o�]Q�֗t)5�&��fho-<�u@��أ?�ǜ�CRk�6�u�{
����!_|�Iv`j�m���� �p_�P�*0���>�hó���Ĕ���!.j~�c�k�S��s>k��_{/���?_�*�PJ�ˇ�P���R%� %!�~~c���;�`cܼk �QǄJ�/G�9ŧ�ݧ������V��5e��,���az鏦H��I[��kIo^d]�(�
]B�}jL��O?\��F�R�����3��N���P��_�A � 'Zn%���S���pqU����k?F!���RQ[�pBᙈ�&Ѕ�)�������(˿U�R9-^dH�֏x��I������y5�����3ʥ7~���xŮ�i������U)s B�p(�=�Y��Vras/]_� �Y�HU9-S�����0�dA���U���h)�g��j�78����ѥ%l����j.�P&X��(x]pj�֤�WtRx/t~��=֡cR�nC]<r`�"���y�{�Nh���S��,&�u�`v�:���%3F�L[��n����r�����=�U;�������u���m��|�%ߒ��a@'}&u�qڠx�#H<�Y�R�pY`�C���a{��&�~Z,�u���b?�D�Յw�jѮ��7�m"{A��%�@��e�Չ};8QL�Z��KM�8'Y�J��l=8���� k��H]�.h#. �_�^V� SV`�WYDv����P�_��IM䑶�G�Մ����{�:�$��Tq�s�E'>6��dm�F'����y_�m�٘�2p4�ǎ��9�D{a�z��~����1�Kv�E8�&�#�Θ��˹"h�%����l��X.��j:�@n� AJmѮ12պ�ѡ~)�,�¿5Hn"�n����~�;��a���[�x�p:�6��a�R`R���غ���|a�b|c_r���,���kC^��2C`B{��	�:� ����&��T�Z
f��Ob�QM�����Z�z��n��ʅI�V�j*\�v�v�V�a�ω��N.`����%����vD�!e�2�? c����"�}�w1�0wG%� �9¦}�6��Ei��M��5M=�^'��l���tn��[���G�y����S�.-P���>�d}xb�u�_�G{Mtq���b&�\S*�f��g����jи�*3���A�k�xl`*UAs,�ͻ�v�1�k�v��v���[�\�sQL�bU B+�_��m��Y�/����(ˢYtv�����)ӱ؀�^��ȃ$�c�{k}�8G��-��%�M���-\;�6�;����cI
�l����#r�8Ⱥ~fh��O�`��I�w_�^�"![�����g4�Yb �n�z>`���GC��LY�s��q�v�м��u���5M;	�"xXH�uB�_�5���J����38������$߆
ٲ_bw�@�A�A����{���Ã�>7�FA-x>���7G�N�����P��k���� 5���g���/$�K��W�8y�sԐ�b�(��4bS�Y�4��p�$��ː*D�"=yp��-Zs+����A!�����'��`M!З� (ZOhuޙ^I �W삘� �XBo��u����7�ҷ)�)�5��p�2I���m��3Y oá�t�بȄ10��q68�x�����+�RYW�� #? ����1���?�3m�=�)'&V�%rkM�O��r��a��P���̔�7T�#��Hf4}IAo8����A��{���Ҹ�ч��6JD�����&:gRn��936ӏ��Ga�Da�3��='��Ƴ���K5٢�s���&RZ��,B��#�)�z|���S�ň2�!	��E�xr/��<��x$�b���J%��o��SW��\���n�
e}�*�p���|sIJa���/���Or1����^E��$A����AG��i����i�j�4����=y8s�+�b�`��ԪOA�5k4J����vq.jF(O��#�%���������<�t��6����5�X�A��B?7ɴ��0�s���80�!�:����&�q�;��	p޼�K��)n�h��:�ds�:!H�A���p���`z�v:������6[�$&֨�ۯޗŐI��N�p���#���:�}�[��4k�bP;��{�i�h_��,2���g�^1���?����L�����>z�D��:$0/ ��$�>���r�|�M-����ٜ��A���þk�3bx찢a� 屶�s&G�J?�3䃌�Jܴn��*v�^��j��-�	��ag��b���"��2N�	Q��#�l>�WDM6���\�8�\3���-e� 2�'�ɉ�u���Ӧ�kLy�R���:��ߖ;�͊}a�:o�����+!��l�9"J����v�Z%_Q����|Z��1]9��{�cI�7�v��s�X�1������@$6�x;�kq��(��I��*;T���^=I|����b�8H��f4����i�!�!�!nQ�1�+u٠&썂���(4���;�i�1m��Pޛ0�`l��JvƧK�p�����2[�~�S�p���AѾrl�a��j+ٰR/���1�.��u���(r��rnz���j
�����'��ɩ����<��~+���)̈����S墫������(���<���f���V��"���_�!�1,4���RP."{z ����f<H��	��v���xup�Z_�~� ���UT%GT	�<��)���c*���Lھ%d�/8X�A�b�2���=�3n}��Z�dO@tL#*�Pk��@�- _h�i����.a� �f󳙐���)����g�GU=����R!� �@�vې0f���cNQ��H$l2�^�� ��|��T��`�� �{i�@�2h�z����_=_����$��N�G��&Tƻ�����T<�9�b޻���P�����2(.��[��q #���0¯#�-�g�f�hy��Ң��ҏ!������	���̼:|*)���	i._pv��y!:�?��{��줇0�7��^˳�}��ږo�*��&ԇM�kC��w�2�ܩ9n��+����J���[��?p�Z�F��lХ�D��lK�aד;����_8=��+̸�B�@��
����5������*!Ŭ� �<�ʁ7.r`\�$0?��<��OXH�?�sX?a�(`��I��߱n{P�w'��M������:&�H�b[닿j�Y�	���y�X�"'qR�O���)�D����T�Fo=9�?�pit�!v��Z����<ƚ2���#�I�	�2c�.	R��� ��f��������ːo��D;i��lA7&�3^/D�c�s�$��C� o�u&zle���h��0B��̀�Sn���-pػHu�*O%ض;���1,Ut3��>��!j�N���RB���4ꂪ�U7O���@���t�BP��l����^�Q��1eq~�V,������j�l=a���,p(m��^Al7W}p���Nz���<�_4�<�I�1���݅��\"N`��x�Bn�\��C��W`�����(Z=:�Zpp������x�*�e{�˂�iA�Մ���U(�:G������B�V�.�������Z;Q�I*�v�mP��o�z�g�J&����,�����rϼ�f�