XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���wSP�O4��d�q�vt�*��R�P6
��x0Mȏ<���J�ձ��=7��ے�Dn!!�Ϸ�W���Ҍ�v��\L4�y��<������s�g�	S���eU� 3�ګꅯ���U�zRЉ���?_a-_A���"S@���6��ߤ�d��ʧ{,^�8�0o�%)����wB���˴���L�'�T�R6}���� rWpx�d�ZY^,��8s<ih�bް��
��_���y��ѷ���sR�_Q`,��Gw�l��d�a3W�M�j�g֎}*Q�}y�����#��8�gdM�œ'�(d_��CN�E�.E�#�[R�ը��)yl �Ț=�b��C;i�����^�8ŀ�J��z\l�~�74y� ;nOȦ�ߡ��s�@��v�2�w�g���'g��>Ƕ������H�_J�M_�K^a<ڷ���+�WD�v�b�3D�$`����b-۫�g��]H�&ex_�b���A7&�<�7�����yEtS�\O��'Y<px������üW����B�f�+r���c��1#��D�Q0�Xz���tX�Oc���� 	����Q�d�C���k�HΌ����u���E�C�V�c�9g�V�O��\��X��t|@"���������#`T�������S���VyЈ�^ɤY>Iڟ���F��e_�+\��gT8Tsg�.ԽH�)6�e��X��T34~��^�t��p�tg,Zi}6��w��Ei� ]�?)XlxVHYEB    6346    1790JCq���F��<7͜��5�&A.��!��� ��	m�sKY�Eez�!`��D��x_-��_���#^7�D3Q�1��~��6�u1ҊzWE��i"�����Z�ӈ�a�y3�d�c����ڣz�������Z���ZL��ׄ}�\��VF�,�.v�gx�>���z%,\�/|��\�P%lU�c�����R��w�ƈc+�\�㹱�Y�����İ2�b�|�`�B����0V<�Ӓ%1�~~����RʃZ�aQ9V��&��4��o�.��Bp�6)���@փ�O'�7���$��E�8��m��ޫd�h�^��БjRّ�7�.�����������*P��q*5�IQ�ۗ=��kڗ�w���1]G4��Á��̖��T��������tE�&A|%7��ڸ���x�no�Y�ŀ�����5��������8K�r'b)�_@���d��eƜ����י�)���X������Fn�o�k6��"$�2d��9R2~���^���G�n�z�%i�C�U�7m�v_�����P���AɅ�O��z�S�K7�KB�P��s�:�}����b��'�@W��Ռ^������Y9�P�&6 �#���E��_ed�^ƸZ��Xw+f�����R�y��D!��s��w���en)��r�ퟑ�p��ۃ�48��n��v�N�(�.�c��(A�:#�3Cd�	�S�ެ@i��+9B��N���{���pF�ed4��+ԙ0�,�"؎�P�5
��g��X�k`$�cOع�E���W\��V�G�`j��c,�'�)�Fmϐmч��n����F
d�[����,������̰QzLv��e6V��/
4�y�c��5K�H���_������˓;�/���>���/ѸI��h�������IF�Exօ�d�s��+�_��d�A���lzKu���X��xd��]`vo#"�f��$��6;N�wp�Y0��%�&���)��U���d����m�}���b�h�E��Kzݽ���i�29x�;!:�XK�W��ŀ�Ke��~؁G�͘�Dw��=I9t
@)`��ƙ��*�_�TKK�%�:��C#�&8�R���-�Iqݟ����Nu1J[�����
����nr��Q~�]Rپ��Ί�}�C:� X�)�Hz�NN�Z�#D��}`_pC�. �<��=x�����E6!��lB��6Q=��Z��ю9��c�NQT�	�es=�D�Sη�(�ji�F-�l5�(�~��Tq���?H4�_\�.ؠ�ZR}�XJ6�h�ӡ���f��'b���3=	n��5�h�t~���X���(��6�Γ���\�=cţ^�WW�+�Х#w�3>�nAcE�"4E&L���ɺ��i�W��V��}�z�GQ4%ظΪ����)΢>]!Řx�>$]�~�'�Hr0x4��5�]��;*}���	�[%�����WP7�(��"��])�(ڙl�E�t+~��Y�>Z%�=2{ƌynMRx��r�o���h� �kHf���I���FPD32�KS!����1���[W��z��+�Z���.��b���<�2�U]J+�"���?��E��MP��4�)��q�#����
)�C�i�a��h�Y����s��e{'?"�K��(=����Ѯ�n�CY��G&{o���WF��<3�	��0�}= ��2�yK���ã6�3S��X�١2�ݛ�xiuH��M�7�#_ָIEڃ�t��P3��ɑ��
�YA��c��E)�C��F�.5�`2ޙ��Kw��\��FQ��RB,�̹[Vh	O�[�pa���ٻ1�ӽ�k4\m�;o);�bDP�?F�ɬ��7ո��}�]����PD�OR��Ec�<~,�)�H� ��O�ɉMb͂%d���}p���\c?�(:$�3�B����1q7�Q�̄�JU"=⊓���'��$yVKW�=���\Ϙ�Oբf�߆���NN�F�F�v=Mٷ��R�Ԁ��PN�c�\���V��Ӟ'�����S~���D�I�hs5�JJ��F"�����
�B� ���P� n|��@Dgu
5��Ȼ�}G��<�:C�~_K�۽��`�t����J���
x`R�MZ"�F줨n����6W��/g.�~���Vr,�2`�|]�/T�t�
x��p�^�)g�7��\|��4�Ȓ4��E�Y�v�%I�va���E~|Tf�5�(�x�̊��"nS���2��K�rD�hL�~���nB��=�4�A��/��K�#s'������<�9^k.��6S��Ӄ!�6)�[�d�����~X��Vny}��.�)g"i���X�fᴉ.k� ݓDנ8�6���@�d��߄,7���y�=8آ|vQ�A�/��X������L�RI,�3Z�I��_���N+8�#�g?oG��"_��hj����&T��)�{T�?ݡP���D�qpj,�Z@;ވh^�D�� ZNb��,M,7����ɡѠ�����?���k�ChK5�O�o�,+ �/6�gl�#5��)�=�o�� %F����
Be#'�mi�u�N�np�ȯ�@��q�8f۸�6��ѳ�!�IsH���6;��oMSwCYQ ���B+4�́v}ƪ!z{~�K�7:�
����(��m��d{�U�� �qK�w�0�hJ=e���#�o1%���=t
�3$Q�4������%M�]w��_Q��	<'S�ݞ-c���F������8NX�:u��VԀ��r��mB+�0�×�n�͢U�W0$c�G�GI8E,s]1���GET"�W�T�o��0<%�Xq�&����d[LJ�����l�ԸK����ƃQ����m��Z��(�KC�`��j'U�S5��"\X0�gp��Pr�>�Y`\}V������4�{@�F��ST����M��$���x�=Ď� 6��o�Ngb�8wtz���Nܓ����j�@k7N�=�F!7���,�m(��r���4ڒ�R��xz"
�sИ��f��S���l���n�4R�����t;z9�HB��v���uS�Zx�#v�mm+b�'F���ë8�Ġ�Y�2��7���f����ϱWW��\�'YM�CC����+����\2�����ߘ��7 ��CԵn0�ˁ�eŇ�G��A ��*����<�XE5!Y��5Wo�?At�\�n E�J��'���4��U�"?�$��W�Y�a�q�,�}�_H�	���P�4�z��3�U�I����e���T�E��d��O�,��6�x�ѧSnc"R��p�ծ&��"y2�å����^�~\(�~��$?����n�;�jfe`�榡��Aa^eN��e�۳駒���t���������Mj��8:��ʓ��U�4�o��j�K�LoQ��PMm��H���>��ɴ7����>�$�[M���Drdڝ���Jl����?e��\���b���ӻ���y�󿚗�#O��ˊ��0�.G8��S����%���<� 	�Z������ �v��*>=�Ƚ�.�2u#:�yyTΚ�D<)�
~�㥹}��D��������[��h�A��N7s\GVD��ڢ���+�D:��Ѵ����eܜ�;:I7 ���X(��ě�z�����U���օ�/+��9{-N?u���I
�޾�g���ၠ��fA>�z2w��a�]��K"�V#ˌܴ#QLv�9����A@�Z��3F!��|����[��^�䅬f̣�P/l��{N{q@�^�""N��K�re$Y\e�ݐ��A�F�ŗ��׽��g"�<lc�%5SK)�l�;����)�{v������?v���R�j�#��%�2���{�ү&��Ԫ��^	S�皅�%���ރ�y�|NN���X�U�)R�L�iX�����w��Nt�	9zU����!�R�;x�"U�@t�	�i���
[�=���i�Y�7�I���י=���v^n
Ւ�_&�|´�W��M3Tպ�e	��3�,��DM��i��5_�u]�4y:�/j�!E0�@M6���~+.Yl��&L�07�[�E�x��Zy"Θ�w�[̦O��|i��c����6���ݳ�lb����y�}���r�[���tbӧ��6�eG.oJ
��~':��Œ��~3��9%	�r���j��w]��i���ɬ�G�^F�3�	xi{#�<!A�x��SK���To =2ۺ���:	D?o5s��e����{�(���gf"�;�\��9�+u2f�R�DA!:����3��J�	��]�$�'�LM�_��/ˠnMS�E��ьA���K���G���Tف��-uvR9I� ΀m�@��ŤJ�4�"ܺ�V�J�z�{GF�u��!���t�1Iy����wW����)wJ���qk����F��~����t��D�f����I,D�\P�������ײ@^x���Wn]�?���(�ɼ��Z��E��8) ��	[����!_���ͨR�v4���8��m�_�`�7�I�;ըG�/������ⴁg�)X/��j��k�\@Le�_eBO�5
�X�a�=6����o���<��y�_V�MP�ӗ�%���/5�Qm����N�Z#ٰ���g_i��$t����,�c�_1d�|{}�F�D��}�V�%׌=�&���y�L"�(�:�5��׭\����� ��[f�-��gϸ�m�PJ
N�a%km��D��:�`�=�FRWX�,��<�n^n<�e��m�_]p�Ky��?����/��έ��F�t��z/mߗ#u�h[ޞ[����Q�J?z�ǵ����^�y�7/鄖�z��]2����kG��߿���R�@Pu�R~f�W��D	��%��<�%�p�&/Ǆ[y�����1�"�Ş��Ro��X������D�n��&���K��
�ֺ{����Xӗ����cs��M����	�u8N�V̹k��͞�`����C@j��WH0y+N��@�|�TSiz�Uۣ%)U�M�U��b2�D~���.l��}Bo臺���~�Zy����3��;�����xY�l����2<��t�P�FT7�4�$ƍ]&���'E(j��n�S��rqm��g��ʿH#<��X��X��{o~�sR�S���-G����`��6X�M !Iz�B>\[?Y�@m�.�P=5������/�m� ��7�WT(Kxv�0�L藀6�D�q~��u�cI��*o������ƚ\���;�-��gx�49OJ�w+���4�ϣ-& �Q��oM!bN{-�#龷�#����}Q���Ӌ^�P�n;�����v��c0�Ga��������7��;��,g��b��n؎���Йm�[�٨��򒒉�K"�, �l��ə�$�n}Щj��ȳo����lB��Jg��I��M=٥])k�&C���Mr��ݡ�(�,s�3.�������la�J�:/k��W*��מ0�=B�������L0"����pE�c���L��ܒon�py�(��'�bR���M�
)&�2�t*�u��c���/@s]�^����ab;
�&��*��P��ť���@�&���'�CC}Ro��I�\��p�(����bC)�a��;�I$���$k��kg��U��\�벫�"�R��@�*�0f!s�G���5���Oe9�\����cqEXZP�cޞatđPvĉ '��X!p�,cm���J�6�y��tw�����+��Ŕ�_U���k՚z|Dp�e����[��s]��o���G9� �#"9�W��=��&�$�zr����n�K�GB#�²{�X2��OA�u9՚��eg)�Z���"�@�X�V(�ؚ"�r���_C)BN�������)i��INd���¤�j�d>}���1���Oc�^7P~��	Ism63i��GFh���S�^��&�w`-���R-�f��!���O?��5Hi���`�;J�7x�� 9	����u��Bm�;�[�͏�+j/��R��	���$��ү�Y��;pk��