XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ܤi��l�
��5;�����<iye1M`�|X+���ߴߨ$�uM`����W�{*B��νG`�G���D�Vacd�gU�G$L�\�j{�������0��28;���H�f	��%Ff��G�rMG��t}����܏Վ�	�I�=�5cd�3�s��V���wW��:|z-���<|��Y��;F; �w'��S�z��}O�����4����b޹�[?W�\�rM�s�U��(��B<m(R9�]�Џ�,�Zt-Vs�̳���g�����+>5~f������Z��0�=t�ju��(��-�,E��������_g«Nb%�l(�~f�;�K�����}rI+ٛ��W�r0`P����L
@�nw9��Ȇ,�`K;��*	�(���Y�9�*vm���UkHnh�U���[Ƨ;����h�9�͑]�%[��7QvWFq�1���X6�� ��0�`�C:��P�¨��L]"�yӛ���O9s��Qua��!P/Ҏ�L'^�h� ��0�IFͽk3A��,�ۡ��4���fG���zSіR���L��8Ϣ��c�Il9a�ɒ1�\w�0���[�ޝ8�ߺ�؄���'&��@���r�4�Ƶ~+��K����@���ׅ��R {g3C���EC�m[�<���b̥^�������h#".W&c0�0߅�|C$�eW�RQ���]���;��ӫq�^��y���jl�@�􁯥P=`8!_&���&h��+��yFI��hb�>m	�XlxVHYEB    a037    1fe0���O��|;}\6�)���,xѠ��ĝ�RDm'�0�nd��ﷄ���`��,����AR�.N�zm�vGa�mק>g�ޜ[(�9��0�����C䃘�L'DF��le�YC��[��<|8���j޷M�k�BM4R&�8��vP�@�{ڡ�i#�P�>�o��M�㏔�o��w��c?m�F~Dd��
(����	HC���d�iƪ%&�/�ֳ[�%�������)gQ�v�5�îak+�d_��,t�iHi�ϖM����3 ,��J��c��^����n�j�5�� ��+[�;M�F�ʰvB&+�CB��1�����l�a��z��a�hTY������Z]�a ���z��7���������ʎ�GTag�8��0s�蒠�%�`2�j�T�uX�9��e�R����X��V����h��ʭ���{�w�lw�5�`�q��/�T�#f����'�u����0��齝յ�F��;�j�Y( U͉4��.��$�Qe]�_�:i�r�p��<N�ip�3JN
�E�8���Ĺ���M�1}�����S�n,���$�F��j��Cs��g��@�刲σ��e����d|�
Bk'���),|��I%9�B�ř��tj)���3E��r%�v��h "1w0���Q�2��UP'o(���!��}}��@ڙ/Z~<�Wk�&B��ƕ�ˤ^�%C�K�s
?�3�%��ƪ[܌�p�c}>��N��N���I2��=��B��=jj�=�s�K+�2�2�|��X�V=!s3�4��EL9E����jP+I����^1+l*�7>�g��}�i��O�1 Z[d.n�N�-�?a�)D�W�l�\�i���~���Y�E@ٱEJ����5 ��W#T>��)H�mo�@��|>{�n�Uy��\\�l���+[��	m�����*���'��|d���/�LV�o�{f��e\N,��]���r��µ��	�X>ےN	oɒө$��-ʔ�۹ ���`��,�s���F��P�@��=�vM����yƮ&�E����W�Iy!���@�'"��z�_+#ub|+g�B��R�5%h�]6X&<��E?Kc�pE�L[�(�N2�����k���p�����X���=98�/'���c�k��zً.��L�\f���&�������������ˑT�~ӧ�6��L�[���݋8�Hx�eǭd�Qh�y�[���I���gd<By-"`�'��8חw�����*=.��{��.cЂ$`�%^
��?�~�s
7��m�ܷr{���rck,�F�0���h$������6N�'9lѿ��r[\����<�U����e�zXk�^��s��N���J>hκ����	Gtӎ���ҳ�x�9j�9 ��g�-�B6`��s�X��^I.d �� a�����N���z�2��[���o�������z�`�������^�ɝ ��cL�g��=`X]��\vEaUX"������
:\R=��>����af���-
ʸ��n:�t��[�x}�3�Y)��K�tgY��K�|sf�����-�֏^����bb�K���s�rKb��a�wm#�֬�_$Ǉ��C�^���2 N��Z9�*�)�l���p$�c�]��I�s��J���GIȅ��f0�`~'����/G�랎A�*	|ݣ��Z���Թc?�W�_��%��T���� *�7]���J�O��($������e��W���y^��r#>�8�s4� ��?}���7}��%;�+h>S�} �DbJr:,cT'�)�@�A���1���X��\�xZ��
k@@I� ��������8�egK?��I`K\�W�ƙ�׸����R��^�;S��`T[��LO�á#A#FU�"4H��s͈\��A�e0����1L� �Q�O���^�砡�'��1U�2mX)"���j��\2}q�ȍa�0������Q�>ht������Eʈ���i��/g��r�n3cjd�ȿ�1s��0=����O?_����Y���/Ҁm���o����	�8��}.���'�n�O�əC��L��+4�@�y�vm7��D�aq��[�{�`)����-�#+@�0b�hC��+�Z
��g�`�q�"��G�8��J�:0�P�׉�F�A��:�&@z��~�ᑛ�r��>�7���#ǟ�ο�h�^XD��v~t�R�&��>�kᗒ����ISFMa#"�k6nI7�#�$�^���*��%�IJ��p��M��kK_����=�	��z��r$��pS������SFZqAT�3�Ն��f�g������{�(R�OA�dE�S�(\����|�57no�嘒�r%���گ[����gI/�T?�o��j���=
�~��Tұ8L�{	f� �$+uZ���>w�Kž��{���� ��@|0=[���XX$��U �
e \�//�����?�,��v���X��:π�8^>ުn�� �������Q�N�	�#��t4Y�7,e]���l�=��>-���.��+��Ӿ"����'�������ӟ��!���+�4M9�{��k��g�	ʾN6fGe��RD%?d� �]�r�K�ps�̑�멊R�����,�Sr>)�,�ۂ�|jAQT�(e�{)�C�T�Cc��3�O^����_�V��j+@�#���Qvw�N>帊98T�dt��I�Z3�q��^�XG����$����/����
��9m���6���w�����H-��i�N����� L��C���^���ԖR��; ��"�a������ϔ�u�7��5��ߥ�j"�%�NUƿ�N��Δʈ���PM� Ժu��n'�{��қr*�S�yt�Xo����G����aq��eG��G�t�-(�s1L���nW!^Դ��;Z�iN��	���k��s�H��Ws.�b�{n6��H=�m �]r�Tg��^���F���A!�(Z�)<���Q>�2x��\b�)B�pFu�"���KC��_�5���lE5_�\��#"n+�������v�84�]c�Kz�Ѻ׽Q[X�A���r�7;�����>TD��00�),�U�ڄ��bUO2����K��0\�;�V��];R��y�d�H�&�{uST$Ĺ8V����2Z�w�o�gOE�%�9�x5X�r�vR�r���+�=`��8?�CoGba��6YZ�>$�$�����|��9��m�Z�ܨ	o����}���z"��L�F,�t��P��>_�2"�d��X3��>�B�\)ޫ��rt�2Ӣ9Z���7�Xy������j�{�i)ڴ��b$��g�B~�h�0��%7t�%�J#�}�j%YA4��?�났X��}[�t&/�Ni��J������<���-�΍?�Dc��=��]������<}`F�eC8�QN�*�9�ؿ�K��r?���ɣ���(�?��m���v�xѹn�/��6��%n����W��[�b4�;�t�co�H*On�O_�r���?��D-��2sǝ}�5��{�.��?tf��{M?�9x��C.pn�j�x*=�̋Y^�۩��w)��~������
�,��¼�
 �G��w5��eC��Y&{y ���<�׌ඊzۺ@8l�}A���h���v@h/�M;��+�����BU=���@��P�d�����vsm��qݿ�>>���)�SiI�Dۨ�cw/Y�*��ީ4�f���1��a�-5M�o�I�uè����U�5(Ed��nJ�P���}U[��	���9�(��;����H�J3�\L�A�'��m:���[������2 22�x.W��×��.�9�pI�J$���A}���S\���4�K9�U����=�2(p�4 �hFl�L�a`ɛez���:�N��FP6#�-�L?ӆ�6����%��Q�J��}��C�k���ݵA���\|�f���2�tH&�ۃԪS?�Q�梏J�S����G��깕����U4�*�Cҥ�����dݛ���'gE��'H��{��xh�cA^.�������C�R`nϜ�� �|��Y�p��^�U'/�]��31�~���qN�-�H�Љ5|�.��#CP�@Fϥ��e�ӝ^o���J���r�+@����>�����2�?(���S�h�cG)�3$�s�?��������͸=�o0DM��K���n��BP�u��c�	�,=2n'n��h�6S]�"������|˿�S��kY��:k���`�Q��$�\�^ �M-������&'���1�f+�~�v��G6�y�7��o�UyE}�Qd��S6�(2Z�ٮ�}��hM�� �᤺����֠�H�q�I+/�dfqM��nZ0�0���_n��{�@b�&I��7>k�]t��(E%mʻ�<�o=z�L?�����՜�A���L��!NBQ�p�X�� �j�D�3�>�`��������r$��g"59��]S�#j&I����w� �|��m�߆��R�]@�����zc>J�N|^e�7���G��A��JJ�	
�WZ��v�os5�?�y$�c�3��:7���B9�	�im�4II|�H��,����1�ax��aDc��{�zj1�3u���g�菎�K|^)7l��ʿ*�X>Z�C� 3�0�<��4r��]1�mJ�Gq2��L�B�\咔tc{�f03�F�ebO^�G���4��\X�9��B�����7��6��HYe�0�8�i���[}js6��A����2>D��"��]�L��}�u� ���c�|���{ 7Y�%�z����2K��o���o����;d���E!9�8PZ��B��~�r������$�)��Z�.�}���|���˒jn�ĩ��I�����YY�K��B���gV!O�%��%I*$�s��}�bl��!�ޖ#���R$\J*��V�k�;Py�W��dX\xj1����1��P�ؖ��-�7 f�������A+��9����V�k�s6��)��Q��UEJ(�#'���M�-�#-H*�K���ooǰ�pb\�W���3_Vv��`l��������$7��2��0�w0�|�Q�,��H������%ݻ�������yĉ�h�7
��MYu�.�R��6��`��m;q��V�&��Ց������FF�+T5�3Z��PG��6�n��&DAU� ��aKb���a�ს��[Yo�q�,���#���k_��˝B�b8Ǥ�DK��	��_�D���>��hD�?G�5�%SDR���h�z��*\�l�B���?��Z��\�v���d5��y�*-J��0& ]3������NK4���9{A�M��<�I����2�-v����f�>?���W�"����aM�Uu�?t}���~�2aj�S�.�X�/�[m�C�jЎ �9^9���I��0����i]����N�.�"��OV��lzJ��Dl^�<�$v�-va�}�|��� a����Cmbm�:Y�#�(�6���n0\�ŭI��G6�$`mF{i�ߟMx��!Ƶ�<L��]ꚪ����~�w6j�ohU��ֈɀ]�>	��*=z�y�S�����aq"0��mO�n��Vɓ֥sL6�F{.r=�/"w'j�&pJ�Yu:������i���q韈ߏ�v�6j���`2z2��O��u���6���Xn�R#��K��]�S���E���N����5�l�$�I��pdT�z�^	P�yل��z6�'F���w�_�2�A�	C�=�]ϓP-A���
͕RRɪY"B��v$�=���_�Vj�T��>#8]�q�j�;���k���!�o̲g`?&�0�z�FG �s�M���lKI8�[�~�<bzC}�����D�	$�,��k�����!�8$�z=��&V38qmy��'���b���k2�P�)�C��[Ī'okf�Y12X@���
�xB��9+�`ca[="W\){�-̹ޔ�;�{�����W�!�/��(���N�ml�Db=�{'F-Ȓٴ8��9��\L��a"e0�t�4�:`E��.ߵ�s��!�HJ.��e�w�cB� |[�����1k��sf�;�'��U�X�v�_ӆBj�ɂ"�އ����;���2��O��hF|������������t�U:T7$4�?�P�f�~�MW�nmзC1�(v�: l��� � �d�z�$M"w��#%9e�n���%""^ƎC��.�$�%���X�fZ\G�k�%�U^�<6G1���/:�w|J�鋱0[�k?��!ؚKe2E�B�&-۫�# �u�u�p.��&��o�@�P�������+�N���vXA�F2�T\dG%4M�F��'C8�7\K�z��Lak%>!�Np��g�	ut��rC����+�A�cJ(; Mv��K�5�x��?� ?�G(.�����;TDJf4�D	���i�˝b�k�Kd���w>#���-.%r^a���D8��Ҟ���
~��$����֓���d}mX��U�"ܚ,��#�=�p��dh��8p���i�kG's5�����5J�[m�Kz���Ek�
z�H���gn|=�#�O��e��GH�u����C_�LVV��4��+����M���7�WQ_���nm?ȭ~�G��5�)$�'#�"F��+h4諄-xf�ޢ�:�ĝ�&E�:@��Kx�h�G ڏ�h��e��ǲ\~'ۊ"�2@xW�?3��4�5��tM��9��˘�bd���)�]W�w�,3 ��cܨ�Dt��7nSD�x�b��Wv��ǂ$;�|w���Dih	�<���@Jۯ��ذ�3ԇ6S�Qd&2�|�l��|$�o��s`��n���W(��.���
�'��w6b,,=N�"/6��?%��EeB��K��=�1�����뿞����"�d(��: q��$��$�B�"dw@T��ɜ�o-ZG��Ӣ�c�ߨY4�)a^�w��|��O�w�;P*���mFVu
u������?�\�3�77��ݲ�NU**J���!�<v��t���'`�!4_z�L�	9���~�8ޢ�ke�֬+�3�<�cV�[ɩ�����R77�Q�V9���t<�����/K��u��I������M�gt����2w����V�l�A��6�3st�[!��J�/9jz�{"mZD8�)*��0�y諭��)�9������͂�K1cH�g`���wgNY,?}�5��� �C��M-ȁL�TƯkkB�W �ɧ~5���dW�A��C�:)U_c@�31_�|��X���\�p�-B}Տ�[&W\������K�N�8o��z��-�.�d5X4ᘑ��f&� b2��:��]��)��C@����
��o��ds8]*�z��fk��q=��VZ�{����3���]	���<
_�S��V����AN�����b��&����?IA�W}g�پ)���"���"��M�J�h�$���[�B,��4,�26�^?Jln�_07�r��n%a!!~�Y�rK�Z ��w��﯌�٨��������	h��Zǜ����M�I�8!����`w� ��l�|��+a��<d����}��)�Y�לLh��e.g���P��y�(��$4�P#��N|����
~�Wd�ͤ��5l ~u�.pc���wz��|��8i9p��ã߄��\86��������{n� x�
�~	�o�;n:��/zjC��{����i.r����� [$�2OzRWxîo�?��-�Vڜ�D��w�0;[0Ag����GP�$ˮ� ���3�|5�Zy&џɖ�0ǔ��w�bq�$Tm��@df�������ۃU�G��5zd�x/�|�0�����Y��6���2��O��H�������o ��ȀOe}�"�����h�c?���y ���2�s6
]������	�'���N[Ŗ�|�L��.