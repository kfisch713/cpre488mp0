XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z�Qd��4���c��l:�V��H�x�bo�.GX�P0*P�P�U��y9a�P'I�E o-��cИ���%�4ju�P{��˓r��m���O�jߙ��m�y��u���Ty��&�oz�MA�4����	?����4gg&z�uns�2R��3�LF���p";�X��K�9����^�s�3٫�Vy�g�Q��iŬ85�������f�)�
e!jV*?܄��S�<���])ו��jGW��G1��w����ƨ[�^����-;�<�p�M_Y�d�]���?�-�T��I
E��ť#*���F��C;$�*�\c�F*�3�
==�jxj!�c7�C*f�pf��p�ʊ�2�W��2����2����uð��W���&$��Pw��|�>���������2m*Wq���,C��ΏE��<�	a�5�7$�n�S��1��:��#��HI{A��_��ЛZ3@��Q�agb�O
A��������ί�w � 5�;��F�>=Ҽb���'�4�k=�7��#UzZ�p��q��Lk4���`��
��� W�Eo�IV˞WH�&�&��/��[Z8`�3E��UQy`�3f��H�k���ǟI9�ǺPM����`����u�-j)���?=s�RǦ(�z�%w�p��K��+��j�dy�C2�r'� ���`�x���T��N����T���|�/۝�~'�ޠIL;�1��{���d�+`��R��� T�ٷ�!w^3��XT��w��2�*�(M�::,=:Ə烹XlxVHYEB    dd8f    2160�i��B8�b�+>?��b6<h�h�p��]�.Ҳ^�	V�)�n�_)���hQ�o� U�N�t�QcVk�>͇2{dя6\1�K�g���ok���3Ы�ꪙM���í� ��T�
����D�:��`ת�6��g�-�����	�xW�`��������$1eY.͕۔B�x)��Fh������d)���fS07� pE���z��vD*�t�)�T<'x��潎�3�M��#K!�g�73҆�!��N��v�?U��:�q��{~hcO�|����w���3�"
D#���Dm~�@��d.i=�jS7�l��J������r�eJ�X,Q�s5n�B,����_�B�F��v�����蚙m6b�9lm���o�!��T@�3m������ĉ��Ґ�ͣ'��Ҥ Ã�E2Ώ�8��Ov��a�9�!'�ԟ�2(�A戇	��w�&-�7 q��g�9Yz�)�����B���!�2nP�h.�[��M���U5r�K7g��6���S�9!1�)���H�N�Ձ�g�R?w>��6m|��Q���Z�M[F��^���?��L�XC54�<hv�X9���:S�\Mu��וYȳ����J=��rY�W"�a@�!WFs�Gv�z9Z.��\������)�P�z=�Zjl^|��^�G�����E#�T�g�,��	��	�9��mu:yyxt�= =}��&4kig����+_]�W��(F���(Hn�W����[X=��~:����v��� aQ.��O�ŕKP���'������l\���N��7'���J�e��2ҷw����Rd��,����k�~�C#�����?�L��*�A�e���o��#��}Ͽ��c�,�_��;���^��^���UK>K�`I�㠍%���Uf���K�¡|�r״R�`QUF���Sو�^cF�C$˟H�F����)ȉuAV�̷99#��"Y� ���T����/'����=�B�Q'��wp�����ޞ�������'��/^����h*�G�{�i��0
���ç���򨸫�yb�>lǰ���U�.�`b	�wHMP� IJD�Km�
X��{����`� ����A����Q�s�چb9��&�~�XO[�����yhg,m�����W�z�WYY�uS]�q���և>;��N�kI���ȃ�2�dI�$�\�Kx�l���3���d	_d�rQ�mg�>eGk�~���aX]&�	7i�����N_r|���8��5�6^��c�6"`�1 �mBѨk[[Mu�<�/��	��w�����~Ѹ%�$��QGa��7����Pƻm����)���i)A�[f�#@�h����5eב�(�ۮȸ���W�B�HOg��E��K�_Y*�E��XH����T�D����wC�)��N���ô�OYնy�� [�y�|Ѻ\���N::x��Zꛔ�x�Z89>���f��T 9��$��@�:�`���x9���ژ�WJnCO�,=��nm��d�3��tp��@�\�w'o�[���i{������h�h��B��v�d�f���d$w3��p�$��l��c:�d�8�&���D����nfu�!�+.6��	�u�ZR�_�=a���H�$ʴ�#1ʸI������h�͵�:�h����g��s�%f"��Ԯ��Kꚋ�#� O������笏l-چ�q��>�_����DJ	ra����˯����~�*6��|���8�=���?њܕѻ��".1L��:\X�>!���_s�dӒh���cf��׾��H����]w����V�ph�xp��Θ^�fw�Kr�/BF�������eܳ�t���K��sZ�^�������A���W�]du^�ȴF�0�{�j[}��(��5��Q-(��Cq��o78X�:��Mu�4:�[*�JwX��^�[��}A�sӪ?=�?��B)�a��� u�!]�֠���jP��=�� ��ƫ'3i��W�#5�,c���α�ʣ2���*"�k�3���-��M�J���^+����.��/���c���%·�.nV�S���w������2�a=-	Ԧ;����o8/KRiC�/�$U��fEc��������"T�k1����ZTa$��l:8
T<��9��cx�_v��@2D��-�)Ϋ��+�'E��w�g5>�|���i�Yx.?M�\QUe�@jࣥ�M��=��`ZV�~5��o����.��v��Zl����c=�vƲ�<�G�O��f�v�z�4���LG4�ub2�B�UCc��O�� )Ȱ���;bt�;��o�mK"�o�V'�8�Ls� ��X��;��AB��h��8�nb��������k
�땃u��
�$���_#~0����l�x��~��g��6�/u1�$A~�]ҍ�t��5} ��k#��@�p(��>��Q/p�ش:�8�5�v5Oe���1�;��6��Ҵ�N�tS��S4��
�3�݅�o�W��HAB�W�3��>�%C&��J�����X*��Ϛ�g�('�f���l�Q��x��,�̔7��T��)c�봾|�<0���1���z�w<.쇝����_�ǁ��k��U~"��v��I��IaN��y���1�fY]�Xe{Tm
g�}4��:�
���/���;�I��E���aAIl��F�C ������e�9h�g��b��W�uR��r$H*73�z����{쾙q$f��u�9`].��]�j.(�@�g��	&��zů���_�J�J��
�$��7�+����>�,N�OT�T=Xv
�7T7�DÞ9�m�����N5z��2�p�-),q�ivn�@��X�nԱ>��/�[�AfrJ�ɦk�w�8��X���j�C4U^E-����ƍ�.[������
+f��v�x�ʾ\np�]w��[�yw��4}As�8������Y��W�ʂ·�0D���|��1���0,u}[Q��1I���vz�M���'Ӆo�|�IŬY��p�%�L��e�
v����$<r�X�:�)�6���¥� �'?�Ll��}=q+���${A�t1V�ry����ѐ��<�"1����R_i��;^4np=�}��Xe�X�a�a>��*iվ�:4��ع?±�*��j�.ſ������`Y�7^7�3�8V�$��Y�7%k����.��3�g�kNj�[������<��[	A���9c���Y3p�d&/�t�")�ޅ����mgK�ļ/n��;�f&��c��3g�;�������X�������.�(�g��2�Z���z�FZ[\=GN5QVj�c�*E��M�k8(X;�{�ڸ'� �݂/�fk�UM�N'�%0�6~���a+��m%�~:u*~�܁����.s�a?:����/����/�ZΌ9u��UJ�0�Px[(��&�-2\����WR��*�h��9_�U߭˶�=�D�q[����("#���Zq���W���7�B�K�	0l<W��h孳���;0Ĺh5��wg#/�)!�T'����M��%$�>\���q],��)��=�k eR�f|T�Z�E~t*���aT�n�+�g���[�����w����r���<|�h�~��ۋa��sM".L|DI3�޻��.� 	!��	,��>q:�M��J��u�#Z�̿,�e�/�𑥌Zde�{7HE�1�7~$�p��kLK	�1�8��z� fY�\>q,�E�����8������|�;���������N���FxdD�-���ؽ�v,(��dgh�ޯmh�Q�è({����0v;�Z��g�9��85�69���uv���a.��&��n-��]6|��?�7�(l���IO��d_�\`eE����t��a�;<��I}��~Ӡ]�J��8;]�Z1>$lY?^��P(��rr�r˺3�(�Xj��qH�&ci{H�w�.�������'���k(b
�u�0#i�Xix��@�r}�i��;�T�'��W�n$�HP��MQP���Ӓ����_Њ��;M� � V0a��ۈyǷ���l2�؇"Zs)+w�F!���4JQ�ڣ���ꜴK��B�4�;��*��� ��L�n�keM��B/�[��]S���g�p�Я�� ���R��x��Iu�x������Ir�l�7˕��+��ϔ�XD�h-��7�,!�c�JS���_)g�sU��_ k�A��CFNw��unz��pn`�}L^wd����h�1`��Nq2�>��}����ˉh���(ǅ=�ї.�۬�����\i��4�l|HPH,���l}m=u_ �B+�c^�Y�=lR�׳��\p����9�T׶�m�[m���
ks�X5t����74��yW>	𜂆�[��O�gD��UT��?o���������a��Љ݇�h"�ʔn�����U$�D5E��� ũ�f�����@=s��`i�#'D�L�D��P*t�;	�:xޫǡ������C�q��[a����bc��]u\<��Ύ�/#��%I���*�2��"\�#P�lIƇ�D�ns�{Ѣ����͎:P�<ebh*�| ���q��+.i*M�䜼7m��Q��<o�p��Z��Zb��{�/���^��-u,�x�����5�P�y_^-s����u�4�p$�9皊	b�̳?K��|_��+R������>���"iRҶ������ll��@�g�4��wAⅳ(�E�W����>���Y�f�V�Ǐ<��^���zte�&�U�>̇���Hs��������c��Y�n�\̣�ǨK�_�bA�k��~�a��܋3�_`��@��%�2��y�.���:����7�c�X&_��5��o���Q8O5C�G]�KK���j4ZJ�3���O�CA��1Լ�����|�LJ�u�
�H�d���{�S%c'@��4������B摲��'^����|�Y����Y�87�b��`cF���;X����GzkM�Q=��r<�NZ�B�[��df���8���j|��r4w�c+����R6������:���C��Df�-� �T���+�[�G��,�$;��B����1���j$��[ �T�����!rX���U~�-L�bAJ�&�AI����Ԓ!�!#u���F����	�1��M�I�/��W +E|k��V��R?���0[����MI��f.F���猅�����-�� �b�8�|������sK�إ���6���᱙��N$�b��`�?�k����>�wf�T�t�4�o�5�[J�^��zH��O5 p'�s� 3����DxP~\?���Q�I�PA͂�������w࡟U`���*j�K�/�����@�|��	��7\s
XZ8M��?!M�1�	�1�5�Իj\ ����U��=��N; *3��V�f�(biP�؋�^���"��PCE�̗�Q1�xʶ0�cr�2)�+���-z�+�P��3�$H��,���O�]w=y�_K����J���mf�h�m�%���	D�_���s�<�87>���I��Jk#[�E�
���|���E�Ȭ��8yD�Sw���h�V�c�O}=�9<�Ǹ�B�0=���xRPF��;��=�����Š $/�=%Mb��x഻�"<��jgmO�!��cƽ!�3�P�]���0���9�i�L���r��M��_��m���5l׫)b��r����O������g0�AP�p�=�x��x����e�F�uj�6�Wv���&w�xq]��h"�Z�X�Ek�M�0�&z�A�u	-�����`�yf�2J��W�;�f[!:�6�M��76�-;��4h+:� �����0K��;Ë�y�ӷ�Ô�X�W�ro�7=f�8��@��Ei _�M�uD�ޛh�a�������:�iܱH�"��A��m�T��?�uF�H&�����6��	OJ9<��Ԭ�����=��<w��6�V�6��
Sk��V&㠺}�?��%��~^��]��`V7�Ay�^�6v����v���^q��=�m�t�����8�����,�H'�Qy��1����d�r��[D#�f����l�K�2T%G���ئN����A'�ڇ�l��}c��[�
�f����Sq Y���҅��S>D����:l�������`�B�%)i;4%������G���7;&�_�j�l
b�?d��u?����B�p~@7����Z"�Ԕ�W��}��9��0��j ���5�|g1��T G��%�~��^�-�*T��[v�u،�J��+��T-жؓ��s����u��h˭�Ͱ5�e~J��r��H���**<8�=���QSE��e�wF�g(��w��v^��
�qH��׳I�БG����,��~���]�9�D�kٸS�_�Z�3ľ�%�==����f�
�W�'�`i�_ �tc;���`i�St�]�������:/L�$�nT+
L�ՋV�L�,+��+�xS���W|��!�$�kT*z� ��H?�}t��\�����?�Kƞ`?7O�NB��6�pKv��O�8�L�-��͔�Syaz�� ����'2!M����>_�*�mI���!觠a�m�I=���2�j�?z\�>d^�ՙ��F*3�A&����)w�vɅ��H���!������޿[:r��~PLefǮޗ6���p>����5�t�f�*�����DaP4^Q=?�Vb�ɢe��I�^;#?"av�0���N���=m������Q��X3j��Ǔ�c|BM�x�>
�[�}#@OX���B�4����IIߕk�]�1yRuKe��C.��\��!XeR�9v0�N���n������ER��8黐Q1��V�K������:�5�Y�A鍔
n2�tY����a���Br��$�+V���1��3X �&ìR����gkD�nd-s5~� ���$��V]��'�s\1����L� ^l���J>�)�7$�oD�E��C<����TW-ۯ�5�l9��=S!���^��T��@򨳻�gD�m��7 �u�l�������ZFj@��pU�Y�`'=G��I,�ort[/�b���5qI�����9����.86��Hk�u��0�Leo����<W��~�L-�O�\����U�җ��3�Bxx< ��;4q]}F�l%hiw���^�miZ�*�����ը��%9�\䍃Á2��B�b� ��y�ؓ��qz�
�)�dژĚ/�S���$��eߛ��-�\�2������[���ѵ@��Ï����&��C���]e���~�*�eHȗT���VYgD���-�9������Y��A���������@ɉw�yR�,X�i�K��6Q%s�~W�%�R�2����->�MYL�jXK?����4F�_��GgBc�����?�Nv�͞V��g�(_�a�y�v9_�а+$&�zպ]�A!p����Hh�8�?;�r�$�� �,{�����u$��8�]�j �� ��&BĔ��7O}�Qj5�Ga�g��>2����Y	5�{A��3�nl6�*�h��a)��65�����?�>J���jz`7��׻=��ek�O��_�45?��|:�4�W������� x��T�z���l�GH��(;nkv�B8�E�Zț���&��\����'��2����B�Jk)R�U_�a���2�v�ͤ&�ͨ���tU�aA
���j ��μ����m�m���e���}^r{�4-B�ձ����[4Rjs�O<����f�,�����.�[j'����"� ��\{�]C<�;��Q'�SS��I�"���ct��/�C_|����O�\�?2z��䒛L�S1!8�U���O���RAc�|�0W	#�?uJ��HV'���4bl\����܃�]5��_��k�X�N�����>4�1�YU:�8���!�o}ƪcc��
>�� ������;��tփD�����zbmA9�6R���#��b�>Ү��?�X�ϥ��}
s�	Pߠ���/!���,�FL����^s�gu��cTtTm���B�SOɮ)5��W,�ߥ�˞��Ȁ�9X�N<wm��N��#��;;��&[�M<��;I��#?�EKY:�v�����mV��>�F�ͳ���B�d�V���K��ʽl(�PyMt`$���?������ߓ/ ʷ`�<�I<
���?tf�}ћ%2��%���ڴ&�w��IX�MN��.��B�PH8�mkk�1�����u���b�����`�Buu���� '������`���(#�RhY�k@ɹ$,r� �4E?���&�ZǴh.�O���ESC_o��:mܗ%��w&ܷ�+.t{^ӥ�⠔��Bʢ=�E�g3�?�C��z9��T�]!��(vJ���d�~��ҿ��