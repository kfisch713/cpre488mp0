XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����>Qd�J6+
k�^7?�B��+�no�&�H$��_�1ˠRc@v��a�`����/-�����KkD�c���c���qc���~�bJ�"7��d����ս�Ϯx%N�A��C#��z�BR_`�hqQ�z�
9�x���
�A|uuhO�<f��Rcj���ɵw,�,&��;��L%��ɶ�ܝ�������潻�0$kq5�n.0��Қ�9<*ٻ!�]��`}9��ꯈ�o�]ZH���������VP��
������#� �Q���U$������ �|$�#9�w8��; �����Y���b ���R�~Ϡdq7%3�?�/�&/9�+�)��-��~#�E��F"Kѡk+�-����"VBw��n�.">��P���X2�����G�:~N4 o�_�ꐐGp�U��w�kY��G�,3�S,f��[M~�khI��O�<~t"�@z�^�+o]b%�)��u��&8��1��GΩ@v~�϶L�#'+.f�c@�4��A��~��ݪs�[/ng�� D�{^4�5B�p�e�vω�{�Œ�k���)||ۡJ�����!����"_�$��Et����;�L�a�$��0�̂�5w�Q�j�<�����2��%+�� 1aD�5����|����Yd�h�������D�<��@4r�gr���Ѱ�j~��3����ͅh+g�{H�W���N�ݱB`�^	+���.'6.Ęퟜˎ���!R�!w����|v4�c;F �	XlxVHYEB    1853     810�����X�[b<(u���4��[�F1���Żݫ� �����)��Q�[4����%�N]fpys_�,��8���z$|�t��:�^��F�P���B���j�S�JC.ډif�&1�&.�:q"IF��Z}�����S|�Mr��{@�����Yn�%0a�c����Z"Ue�V1 򦸳;�ᥦ^8�?����X�T��٩�#�T֚W09u����8�����_�5�o�T"���V���f˨Y���y�F������ײTB� '(�@��&'��Rw�����rx?��
�7 �9�;)����Y�h,��Bm�O�q�KZIގ��5Yk"H� (����M�;�>�}j#����}0f������7��/*��Vl�D�֫obg�C��Ï+���ʆg�a ��]�����[3�ú�L���Л�O5������]�ЍF�<XF��(_D����*��A[��&�=����<�0�1H��4M�NMl��`���� N5�U<I��F[��DwA���[�_Bщc���,H�)���=�Z����a'�5���ږ �
�О$p�.��.�ȳ7��zzc�H��)�0yk����LT)�f9j��'��fo&�-�Vz~������n녉T��8i^�P�'�d���HT��Ԍ.#���J+�.����X�E���[����IS��
iyTSe�q���Ü�\R3_�yHB'��
��>�-(��ԘM+
���w�%�..�⡙Q���7��j�H�w7.E�hbæ�B���]f@D�ޡk�I�\�Jb�a,�i����~��@��5���6������^U���l�'�X���e�b_>���� ����'t�Z����)��8�TE&�>I�����T���7wo�_'m���F��B����h�D��P���پY9���F�]�r���8ԇQ��y��Ml�#5��dn�j�F?8���u:#"S�M�!�Ⱥ,.�6@�=B�?)1�&�8�̸����t��	��>b�[~]�U�u��Kj�8��z�E��\m7R�Q�EAyʙ/��d1�L��㼻e�r���Rh�z.�|��h3=��<[b(��磴�]m g��$m�>C�-���s��2�����T��?�U���:|����%F_�H�nUiv�m!E��އ?S�pYc����kd*�y,Y4��䯨���L\��m�)H{��?V�ud��x����+�J�ߡ�rl���tT��<�a���/��Ņ�g�B��V�G���|�KH�J�d��<JJq�esS��S	)�ۨ<��������g�H�?�/����Ժ����:���&-'�{����~��K�r�F��F8~ms��d�W��y	`�S\�Z��Hi�E��1�`���D��k/H�!��i}��:��E�ĭ�[��(
 ֡����?�֞l���8g/(ԉ+�ƌ,��<}��\>��fְ���FG�J�L��9tnK�gc_C��3��>�u�~��U�}QտE��r<'5+��0W�nH�k7��3b����N#MX��L�A\=R?_�ЪTԁB�|������:���8v]���ͲSzw�e��$��	>R�bUAT1xus�v��<���sQ:E���9TC�XG�:�b��A�$#y��Ġ\9���}����`�[d�x/j�eC�~�Ĩ��-9��6�7���,�N8dɹ��h�-��DըF��6��#�S/�,L���YIb�9D�(���6V-ae������=q :F"-&��}
l�\��\1�'�7��EP��g���YUT/���@���W���(-*�D��� ^:��?�{��
ߕ��UWvo�z�("��N�1�Ӣ0D�K�)u��*d4��#.�~''��
�p9Y���y.�u1����[1�eTL�Z��;��61R�Y�]v�rZ�n����
?a�|P;�O|2?SI��3ӯ"�X�J�^�&=����z�OU��"��uL��R8f�WJRK����T��҄57J���xr|�C$���}