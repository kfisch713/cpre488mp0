XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���K�af���м�(��q�c:���0e��Y�w��>,&��{j�5����/.{���)1%=
|��Vic�D/����Y�74�����n�)w�uC<皷T\�B┆�_I��e&�Q���XbB�,RR_�������"��\q�'�\��Z�j�;bv�*�����ӷ��ô+�vZ=hk�^��p-Qԙ�t~|n���KRhCUZl�5���/_��#����Ś�3tK�9�ڶK��:h2f�b�=�c���]�U�,KŴ[�?;�'+'��e�~���g:/��HJ�	U��u>=֒zд��TrU}���3��9m�>�w0&>A�=�p�;���p�p��N�VZ=h���j8�S�Q��8��W��ڗ�����5�W��nh�BW�7H^������^��0����E�R�WN�.�bcx�2�[�S��F�d��e���ד)�ᢙ%�SK����6e���L�(c�h՞i��^ӭ�	���$��,\L�h���s��S&]w�t�jlo�`3���R�%W�G�;�]3#�йG؄1
>���>T�����y{�+aݟw���EG �[�&9P��:
{˕q�nw�/�%L=k`�(�}�^�V�!�?���ȓ8x7�	��!��E�d�9� +UZGE8�OĞ*pm�|iVj�{�w\�nW��>x��B�h�~h���.��֙g�q��4�(x,����f#YL�s5��f�=u=��� �O�~���Ik��'XlxVHYEB    1853     810�y��t�li��Ԧz�f��"KXO	|��,lH��.�V�t�l�#7vnoޏ�e}F����=}��ǰ�u΄@r�oI���y�5B���h�����;������Э�l��Z�v!��}p_�w�J�mD�M�J��dYH�M̪S�k#~߲́/!��Hkp��h���W��E`*����ɷ,�v���_����a�zo�ǭz]M�@N��Y\�e��[����o"�횵<�]g:Jj��ßQ�0��N�Zx�!�������)Z���"� ��ri3#�Hyc"�Xsk](Ŷ����7D�f@%!��"<�;��6ѷ%:h6#⋊���^���S��M�	Ό�_L`*���	3�-䴅;�� ���N��!�znk�?��ʍ��r���Ò�Γ���Ip~W���E��Z��&�������tc��J��)�2�#"m8A�H
��-����(�F�Y?U�+0(�m�v(⇱������C+@��ȏ�R��3�J�-����|<��uR��D��y��q��m%���,<���򪴼��d�Qy�q�����D�(��<��	��!P�T� �m��R�ê��߭�f��P�:2��>e6�a�Of�"GPb֮���`2"�� �����t�;�3"�����פ��z��;��2�hS "���Nj����#g~C�bl)ZW��8b��ӑh!�#�ZR"E:W�7.�U�����XVg��I=��h�A.H��hJ���!�_F~c����^I�6�L�#7�w��� :�7Dl���Q�K$sK1Հ3�PD*c7�����1K��Գ�n~��,Z����X����mՔ�o9�r���I�ƒ_�;Iը9"C�60pJ��
H���l�qrW�pn��K��q��uP�(Hl�lY㿁(��2E��3(��!hq�^m�m��@7�g���G�����c}89Va��`(E�5ē��]����}HǨƛ��4�{%�Ch|��B;�`��=3�����!��{��;F́ST�/�,8\�i;n�������ǲkɭ�nM^�i�Q�.�n���%� <��60K��B�ear�{�&��%yKIqӚX���I� �G��[^�o ��Ѹ�i�ɭ�c����<��.��(�܁|¥RyL�<�aH��8j��ۻ��Z_�e����YR&�~`��vȨ�#v�β@NE#x�=;���ȘV�k��ae�U���e�f_b)�x��>���a�.`�o:��z�͊�c^ˤ�_�����mlW3�oXM��n9uO��H�M`1D͔���T{��2�@f���L%��~������Ô0ҿ�};�q8
xQ��ŉk~�p�l�[^�������0N��[�J:�Z�FY�qy@h�#�����[��Q�y�|�<�Ã�ڏ���4]��m��Rj%J�`�9�<,1� D�yu\ED#?��&�3W ��s��%a��V�����i0y��-�X'�2�-��V�Uѐ��+�Vq
2Gi&���>���#�U�{U��@#�H���ޏ=��<;��C���ˏ�V���ۂ����k���%H�����ܲj����N�&B�W1絩��k�4K+�$0��:��e�-4�^�-]C6xv-�B��a��v�����í=�4���k�������<�X���l�H�P \���a8�*�>��(� zU]�½xq ����)�I�w<�%XaP�|B���&�S��¸-���_V'>��L�p�U4Vz3F2����q,q��7���@7���	�k��S����b�2lR��.h8���j�<�S�vSYͧg��%~a���^�n͵÷#��X����x�H�������+2y(�w��>��X^�U��2���ʪ;c�4;��1m�3��as?�����xr��ʨ�N�U�o�A�o���5i�RJ{�'�KK�녝,֛vc�<�Lޭ��E#*�D_�9�ྦ��B��.<{QjͿ>�~H%�F����gZMhس)ikf�sK�2�