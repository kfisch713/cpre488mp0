XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��IxYԢ$/r����W�TlyAi,���iJ�l��)jN�z*(.cP'���w�jplľݫ=rh+d��[2�,�ۉA1T���h6�k�^�]�=��9͊�u�y��쓗�)�+gQ�%�;�mL������Id�ڤ�}��-�0K�)�-;��r۟�g�ǀ$�xt�rq��p��^i�4��l�{�}W��0��[�+�.��WS��t�����|���B�j���Q^\K�G���q��9)e ��:?�8��^�^/(gg�-���0��"����6~�(�K�7q0��%?�jt��0�@�����o�١�.u����v�˹�eƱX�� 9�`��.žlZ
 qlv����Y�րg(��8'��ri�u5W�TXuڼ�g�*H�D#~ez��&�A(�c�gN�7��~ux�!Zaʮ�؄�^��=�����0�x�����\���Ogբ?�J�:8�TaN�3�!��N �O��,��j})�O�A�i޾�"Z� ��<�Ң��+b��>�FO[4�{�w�Vq����fR��Ȭ�C���,�t�����Hc�,�#+���z
�hK��$Y;�gF�Q0����&���N�3>�A�e��(w~�s�/�Rf��K���~rw;y���|_g�ucZV9&���7�k|l�)G���:�_.����	E�{�O�G�����],'�Vēi��%� ��մ	`����(M��\;�3¸��eW�0���}zcG�B��@���j�.�{�}x=3�zP���R�o˼��V0ŗE�f��XlxVHYEB    dd8f    2160Ç�Cf.�{r���
����o��@)��nBH�E1a�@P���	L�*���mxJ��A��0��f��9�O�EX]���D�ƎQ��5䓀Y�٢�g��c��H|�;����媺H��^[��@C�.�2�:ߏ�j�\��J$��������-�
�!��l4y��MIǿt��%�����!{0|��(�0��n�u6��f�e����&{-�����Ț�	a���j.+�H��e�y��_<hPAq�N]XT�����QWBM��l�=��+#E�N��=}�@�*�T��2������l��Q�E&�9�eLe��,��w�*���R5ɖ�䬼�|�R؇��q��5<�c�*M�'���X�#i��LÓ�u�c�p�qT��7R�{1��AA�_����[����D4ʬ�j��3ҋc	�P�C���g*ΕyK� T6�C�V��^}���Z�؊H7ᢓHa� �7c�B<��؊}���ճ����bf�gY��c�<-���A� �K郟i@l/6�{I)��K.�R_f����0�!�E���[�����Ep�f#���u�}�$Deu~4m��y�,���E�d�'�0�S��3h���z�4`�:`\9M��ߜ>��ZK�*&?�]Y,ɼZJ����+Z��ǋ��B:��p<�Țѷ�A������b���G57�ߒ`S��ݜ��� �e�1�I"��`�F	9����ۢ�x��o����nX��+���@YA�`@l�.X?�}��Ɍٽ=�\Ź|�c�Y�ʴ��}�x_-" ������p�Nc�^fy-�;^�'6���3��%:��{6�����}����w��T��h��{��W�>���k�ps����>��*�U��1s\s��ԣǐOX�3�f6�_����#�aFǙ�h�²
��)�NMI&�p[��?�kH1�`;�z-W�C����5�T\�z�9��Ph�[��tޱ�I}���? ���ݩK�g
��MK��GX�.�U`�������P�.�oԑ�-���r"���Gk�1]���lEj��ӿ�h�8�~p��D-������r'AƔ�$˟��%T�F?���ͷ�Ƅ�b;j}����� �E��r��!�����39�A�Е3Q����>���e�G� �ߑ�iU�	���[��
ê�t"U���������v]Pe�E����n6�|�a�/���Y9��tʢ�*�.�Srr�k���r��N5������. 88fb��|4���ս9>8��Q�R �����m��mu�-���Ú��/(����q��X݄F�}h6Ju!.z���=P�������}'�[�̊���V�n��|�ɫu)�sg��3h.0iI�^���u�<�k����}ol�HY��>B7.+�@v��R���,H���Y��bx����P�n�{7]�:�x/�d�\$����Ӓ:%Ԡ�Q��r��Ԟ�P	ܚ'%�w����Lwe2 ju�?��h>�N����z�;5,���DDC^�_�)�̷�,	�+�ܧ��&Sd����,(v'"\������7�b|�\@� .��
-��7-e�j��ڒͫ}y6��P���2��
�V��^���9�;B,��g@�9H��c��.���i�������=K��I��M�[��[&��B����	�i�A����5kr�;궅����\���`=�pc֍V%P��Al�/�/�j�f� it�(�&� �"�%� 6Q\!4l܊��V/�)d���\nB_�<.]\2uDz� }�����l�ʹ��f+W7�_��R�~b��緉P�2�S��6w�w
�! �9�
KK0WS���{�蛧3����o(��T�@�Q�]�e
�_�\���k���MGjh��K]$�]B�8�#B����fX��2u�m��1_'V��
�`F�&?�i��+U�|�}����X��֍b{Z�97-' A\>��S,��7.�'�y�1��	4b�ܞ+F�4ա1�08��:z�B{{e��3�!&�|fi�K�;����G}��4KC�I��G�F����������o�������g<`��X��S\�t���;0���� �sX���(��/L�s��l�"!�='K��H5U
���\��^e� ��O�|�$�:H��0�h��j7���'8X����>V�G�k����;����Nq�_�6���g����I�?J�<X�۾�C���趌�@�:	K��A�Q�L��#��h�K���s�J�-�)�7%��p����u;Y�{;�(Vky�D�pT�̞G��Q0
x߀�0�W	(�r����%f��I�k&)�����A�=A��̰�pW����2�����q��F`��."�Z"J�Sx������@.#�>r�'��a�{��p��u�}�ܮ��3h�`\��gO��+��]���>��l�����!�d�����e��	 ��v�;�V��u3�1�L��>��u���f��b���R���T� �q_��$(O����A�"�^n;y����z�~>���j
#V�0i���kq W|����"��[�b�!�6����	����¹Z�:Ȅ�mW8�W��@�5
=n)k4��Q��Pl��QB���9�� � O�J_k��g�^����O3��.�B�x�����-��U��ImA'ڜ���a���xJ>4α�m��N���O1�@�q���9no����7֤�����I���d�1o_���x�
$%�#�_�����1.6�
��fbE)�p�s�����{&����+!Ϸ��3�cr����	`n�@�|��90wz��}�����b�Ɋ�Xk�Tx�Hߒ�p*��X�A��5�Ю���Y���î���v%��p�!���c'R���J�N�(�E{�S���r��2SE��.5� <2P�VCg{�Wv���ެ ���cq�#E��r�(��ltr�<��l�D��AN��+�ߪ�a�ۊ�o�$����O��i �:����${ɜ`��}�C�;�T��'����Kv�]V���"�o2v�����y�& {L2�9<������T}w<Z�^���SAH|8�����C���9S�A���j�����K�!�=���d<�V�n�t�WV�vy�@ɬ�z��B�RC'흜wZ`�u,_?��k�Ev�u��7͵�|ݴ�?�Rbh_���3I;#x�S�0��O}	��	C����Q�ሥ��0���:��am�Q=�؎�����4E[�����I������n^�,�a	�	�%v�'.�O��S�4���z �M9Ɲ������RccT�LS�kJ�ND�o�飈6��d���s�o[��	?2)��Ƚ��+PR!C��tNKr�~��M����d3��o82�G?`g�}EGD?"*˵�G�KU��eQ&W�Cw��-�+�^�d�d�O��e���_m�E��X1����ކ��r�D���Y��a����j����ȯ�`OX��U5�^=Dz���Ix/|��v
K5V�(�}�]>&��5.��97��M	�X��[��M#��i�˒��N��[5m�Q��۝�ģ��i�l�}ʺBb��mi?�M��vVhTM�i�h��Oz\����9D���Nnb�Զ�����D�����L�5�)���:L�����Q���x�x'˵n�T�U�㬶�BU�O��)�B�&�v[��$,�P�����&�0�vG|qB�nbjЋu�U�������ob�8,�5��?۰����_Ğ�Ra�sM�y�{S�-��g0Iϕ����?�+=n8O����D�Ӷ=�W�JPhjGlj�,k������b\���z�ax�V�8�G�Q(d"	pu^kMIɃ�{6�q��[��~�&CJRb�N(4�h|ǹ�����-<p\O�5a��a|�o��*JWZ��Ш��YZJB����<�yi����7����WY��:̊9�%��d�[ZG�T(�<�Y����}t�bX�'���S�A�Y�k���GZ��k%� ��$�Vy�'�Pl�
��h�6l��	L����`�����2�Ӫ ��^_��U�e1��c�����_�W�ֳ�(y��.�=uU
.BJ�rʑ1EvdK�K��P�NRo�B <��]�U����V��"�T.�kxW���'	ޜs�N�Nw�>+��G!?�<�I3���O6}�	�,��g������t���v�9��;r�@�(\ŋx��;�0��{}��#.t�L�Q$��4����4b@2�U��%��M{]��ūF9-�������$I�^���x�~ԟh2����� 0�Ӕ�M`����/<�/�E�0�~���A� s<=n����B0�x���^P��f�!Ê�"c³1���t�;7�K�߮�}ꬷV)����|%E��r���{�2���`_T{�{$��0��늟1Y����fc��*֛ �q�u�ҙ��DB/�����Q�v����?O��T���T�Y��R�������V��4�6[�Ne��qGs��
�G��o@��ǜ���fEM׿g���!-H�?�i~`!�K�G�P�J������?
υGk3�/	:FS���Ǝ��tr��)�3ot����4&����}����
X�^��^��	_:!��f���X0������?6���2�|8�M��8�%�MÕ�=B���L\ĸ��h9ƶ�^�� N��p瀝��n�h�}��P�Ee���[�k��5U
6���,�����*0
[6eY�w7ҵ3�*������	Ă7����U���@��Q�Zap�2?����n*�P�~I3Q��wz��M��ENA���A��;D}Q;.�����x��'��\R��;�Huh�fUW�?@28�w9ڹ���t��AO5��x�I��X�i�#q_,�v��%j��
%���a6I>t��1�"B�AO�z(ˑWH��c���s��f�˘zyVB��ģj| ���/�Z�I����Mg���07��
o@!��߰���4�^�*r\�8+%�b�),�Dy�M^��MS�H�wU#���w���kP&�ڭMp��\�d.I����k^��(R�x��	�aU�e�M|���������H
��J
�PMNs�H�W��G���J���?4h)ۿ2��?ϫm�����J.�$�^ZY��;�����k�Y!�עy32�Σ&%>%���A(�M����)Uk�yM�@wE�+j�U��/��դ5�>M���涤f7�~�hy*�Q[ǉY_���a��%<	j�;��OE�����٭R�|��L���3�'�/Փq�n=����d{z������(��z[���
�-Cau����N�+H 8�sYW��b�W��M	��=�o9��ܮ�W[�7�8�z�5J�8B _J<��&��Ox��nN��L��a��3Zݮ@��f�6��4�k
5�li��g&MbR��S�	;J�e�V/�ǯ�����r�ɉq+g7��ZX@Pi�%"oz�A�2лB��d���w�|Jf� �M�V>FU�n؎�L|�W	�Ѵ ����3����/,J��77-4z�]�&`ǧU�
����2N/����E��6��3o��6[��j�H�$�nHp�@���=��n�i���.���eTU+m��{c��(�%��)����|Ur4�r����;.�VL*��}�1mJ�{UaL��Cn�ؼN"��`���2���OzVY���$ve�Z�A�;f
r����R��,�,�5�@�z���N���^cD�
��b�>�/���v��
l������Ly�e�^f�p�����H�X�#�'���H�)��L���R]Ȟf��C�!��y�8����~���X��
Ӻ�.�cFM2��U�X0�	����y ?*4�Y�}�lá�y�������\!4���#����I6K���0�>�S�K&k��Mt�P�.Zs�WѺ��Q���<��"����k>I���̻�n����� �Ze����.7^�c�+��;}=Pl�b]|o���E�(����O��kYZV� q�rf�\Qs�Px���y��p�7YiF?���q��ʈ2��Ţ5�h�ƹ�+����<5�v)P�ї�A�ã�/O�o�wsR-��M�ޗp�̡�j��_�9�SN����p�w����B}��PO\�����f�Eᑙ�v�%�Z�l�|Z"tB��`�gݻy��n�x�"�t���P�����v�~d=� �d�3�W:QmngRO���y���& 0���TfO��/7���5VZ?��qҘC��X��@�CR�4�@:�C���64@)�ee(�:F��Ԃ�C��*s��
���v��gLM ����Q�^��A��"S�U<�q�>x	dm�$��ADi�#p�!Qcm�N�C��	����Ś�F�.n��)}��V��AI�|N�Y�;5��(�A���!���y&g>�c��M�^�sǶV��gqg_�'��hK�9�'kr�'c�������A������T��^�_&��!��P���玦Bk�r.�AR	
�������.�ӥ��ؾ�̇r�4W/�_�T^��m����ƃ
ǆ�p˵+*<�X?,g*>.�Rd�A+8{�O�g�ӌ�Ȋ���#��fD4ObOƉw��d�P��>FZ6\aϥ�h[�1C�0z4�I�)Q��޵^��^f;�L��%�)g�sY<��=6��,��r��ۺ�Ǉ/�4Q��W������n�����<,:0�x�b�L�b���!rQ�G����r2&����_"�v%��=,�k���"EU���*�Zj��/]
q�2���~��+PGw�v_�C�ᔩ����$g w�?�,DP��x�����g�/q���������7������.O%�����E�ߦ+G[�g�<�Ѽ1���(1:��`���	���Y��ޭ��H���=��k@��!x>��3NT�˴��'���4$������G�&b�ٵ>���\ZM W�P�И�(d��G�*�tX\���Q����.Q����c<t�j�N4uG#��㧴�=l�I�uK��� � U1F����[-�.�����y�@
�ۏv�Z(tGgu�-]0m5l��>�[z��%�ay$�n�ݕ�	�����K��ϧ\f�Q���K���@��Е���3��}�vg��K G����;��4�[�E	Ԡ1�����3P�����Ԅw�]��1�׳$w}o�0���_ϻUz�e��VW)���������[d��0H��������@�U�N�n�3s���H���S�
�r����D ����>�V�3�%X���Ll��ܷ ���<��r�>U׹�<�}���Nyx���߱��ׯ$�r��.R8�*��`P�z�)�d͇N�l�y_½9����������Tl�J�ȩ$5G�����OV�T2��i�/�>��Br�ԡ�����d4�Oi���v^�Ce��ʹ4�(6oX�r�p%	Ȣ��.��sJ��֊8�>.�)W$�~�*���ZM� >V?�2��Xɘ	�$SL`h�6+셉�>})44 a�  �
lV��s1�3�� �d����Я59��{fU�I�+ �<��Д~;�ĜA+��`�(Oh^(��[�e�y�wϻ�����,����ye��K�5Z�1�vƴ"��S#|������E&vO��A��xUL��Ƃ���q�Bܨ 6��j	6n_	z�_��X�j�`�8�uh;E�=��8��W�)x^EQ���^]X\�ׯ�9��^�a�E Ǎ�߮��W�Y(n��+y������aK�:4_�9_2E��2f�;�²��5f~�TtΒ����W�e���Wj�U�()6�R��k�������L[�&��4����_uy�T�x�d��2��?"�0>Nj+�fL�D�im[V�V���}^"�
,弩7�iTK/���d������x?�@��k�}��k�����v愋�gHmں��?w��sJ�T]�7JEr�i�7�r���$�X�5d�����ã��hb�t!�2�Z������{��8�^�~�`��q�~3�*��`����mݽ��ǉ���u��
ԶF�t[.�ؘu �����^��-�B�/����χKx��Ʌ_#u=�v����[��5/�z�8
�މ;�O�	r�	�N*��9FI��rۻ]��&���Ұ �k�*��.`�z��q��:��YԎ���!�`oT�/��iG�k��icj�H���� pR�a�i��!
]�N�J���qc���^y�}�V��@e`bu�9�_(���n[�Ei����^3��Lw@?͎8�Gq�t�bs����1�vv��E���!!+���a0��%�=ަ�jh�)�#t��b�fW�S�dAX���e,$��Ս|���y�X/���0��������/��[.