XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~����M���o�H�L��y�Y��u	Ԧ��%�?�d�&	�c�+���2t<�R����jƒ1��X�q�R��H�C��a���j���Z&�����6D�F%w�u(q� 9�GQ3��D�m�/{�b�X���֋��]hϜ��9y^FcI�'�b~�����o�k\�
��-�=r��!�èM���3���
g���T�VR+2Rz���>eNmI�}��)���gxT���nj���A�kmG��~���, �ؚp�x�M;y1�|cA>�y��7��a�|W����8��#J�����6�3E�-�IyZ���m�qI]������3��O��P((8헆}u#��`���j4�N�[�qVW'Q�0?����VAٻ�B����1��2V/�1o�b^�K� �
����Ce����_ ր�%�2��[-��l�E��Ҡ�aty�а���)���WG1n�u�����c�H'tyL���h�:\	�>&*m��լ��"�ȅs� T�%�� N^�o�n��;Q�H"���"�^4y�KZ�d����O�S��٭��,M�A-��5)1��`�sD�|�H���u�P;�Lg�[|�n���1%蛜/��8h����̳�v V��o�| )����y�%����r$�����-�����;���"$�I=K�#�f��5�1d���B���K�.)8o�`*��bz��d %���K ok3ї�e۴�Î0�^}Ji�5
��gE�S�K�4����Y��G����g�B��XlxVHYEB    42ae    1110UM�m�����p�g�m��'md(7�`�G�I���?�E����d�	��0@g
��l���Z�q����a����C� Q�t�^G?]i]؉˒�|�]tۆ��z����0��5�C��r[�!�h�1(�$Y�X}��X5{u���awҟ.�4���zޝU9̷2��	׵����ˍ�6��]��C�i�R2�Ϊ�r:����#A��&_�C!��X�c"ՇB8jLW�--j�������^��`�0\]���?y�[�#+�'���%���5m7���E��5��KHn�1�����|�M骈Ŀ�<�Y7��{v����|�C	l���߸\�pJS��Y�L@��p�W%�N���^�*��U�9�q��n�u S�,S%�sUN����G1��G���Iݒ�0������kɱ���Y�	��[4rL���y�/d��}:�tӜ�������l��7bp4�x��]�"��i�j�
��#���${:��.��1�o�DNs2�.0���і�[�F�FT�{���3=VX��t�����[�6��t��Xd�!k���!kAbW6Ll�����eY��RW^���D����<��[Y���l�S4��)����y)G����zj�_�R}����M���V�O���>UP����i�^�ӥ��ym��n���|��ng��z�(����;V��n�q������R�Ū{�	��A0
�cqҿث_�ձa�w�S�_��!���¥b��K�]X�����&��6;r��>����j�;�b�u�-bx�>��m��$H��BjˇF����%_�6ɛϮ��Q�\|�6Jb*X��:�c��W?�N�^�pF�Z���,��&c��4�2-°�TE�[���X�͞��g.�.dΧ�-�2t���/ %ߒ>����bV��'��b���>�������S��C��8�a?q@���-�X{�>v,�\�엎�3T^ 4�e溷�[
��̛��HJE6�{��ΔH���A)�y�a�qs���$o�e8���]s=�μ���<~e�ϸ���$$��1��p������A��t4	��#H���2�6����D�֐�����*�	U	���f�=�DSp3����ܫ<�KT�}ٟ:��pb�f58�@��0��j\�գ.b����`#��K���t���m-@�8�">�A�/q�y�!��ߑ�&�Ff�c�"�����Z�RK�����oM���CT�^q��}v���ɸ4F��dK�{-�S�<J�9u}_lYX�Z�D�P4�SĮ;��$BH�;�(�C�z(]�+�=���qRCѕR�Nl�@���	|�޿o�ԳY��r-�ހ5UZ��A%[��W�v��jD��Mc�Ϳ�*������ݼ�!hِ[��*�]�I�&�������r�Z(��"\��ֵjW���Y����"ŀ�bf����;�5����H���G��D6�hb�Q�0��G�I���oz���Q�	�]0�J�I�ǆ�6�XOI�D�$&[�E�c^��/�k�-��u�S��4��?!����&�?B֒�/����bE�H��XT�6��5I^�n�}��a�
�����S�pf_�[��d�=�>el�$+�8?�5���S�xJ�)'Yk�7\�V�Y�NH�d��F��'���b�ϧqq7���|$i�T�ŪNsC�|��BF}��#n�9I��DQ(6<�;RĢ�l�4����o�s�i7:?�=E(�ɹιѿ1ĝ�D2Se��@�dzֺ+"C��D�V�.� �r�I�K]��|��=�3��:�U���u[�P6s�-!�E1��'�0�u�ل�ǚ���:YK/�����l@-S�ν�|)�hB�e2zT)�`P����{�ś�,821�]T�.�!�p�M�&19��7Ԯ�����HD�Z+偣��b�ZZ_ƙ��k��ɇL��7�c��	�5��a\�T���T ̜w��?l���*�02ju���0c��h�UcDM���>Ｈ8��7����mm��ҹv:�р�6��_�g^u�����}�`����`�Gp����POVN$�}U���gژ:�8�A�T j<�y�VG�����s+�s?N��zL��w� �9���8`�"*6�k�݇�ط���U�.\j! Z�)Ȋ逞���P.�U%5��@GI�_!ӆ��7��9dY���$9b^"	��H.��N�F϶Ƽ<�����V�i"٠4�0-|��kj��]��bg]:��)6:/�΅,JN鮌%#�&��,��ӂ6���āqS�P�h��݌��Z�+��X�Fӱ�����=��̒-4A�g�v�]��hc���3�1	O�>Sv�4;Q��چ�N���<�$�K%=��L�������){4f�a�#��~
�J��F�RUdkB��8T��%�G�alg2t�T�_f��ZU'��XT��V~�3`9��u(�.�,SB�
�q��ޢ�az�R�!�ɑ�[ޑ����uw7M�X�Qh���ec��`��A/(Y?���'%��sIE}8̗7�v�n���P'�r��q�[t|�x
�G�|��;�{��BAQj$�PcE�LO�P�34,�%��dq[�x	뽸[
c��lS����#�e��C�;���kb��u�L���@�ڐ��9M��P�p���@�Ǽ�\��{�	��03��G &��@/%C�萨�!�C[�����)Đv$b�"�R��H��۾�Ѵ��dnF�R���Ci�(n���}���Te������eӏ����
��RM��۞��,/���������U<��fi���I��]�G 8�!�6}k},�@���ƶ����k��@B�G�+�
��7C�cp莠y��|�!@�E����~FCၛJ��bg�坕b�am#d�f��-��\�Tw'<}1`!�͆j��ﾉ!��5h�iXCv �R�4כ�ɫ��<����z����z�u��g����¾�b��D�@���;��ŀ����2�W��R��̎"Is�)�^�M��a6�V����Kr�����d�Žm�����.B�K?���d����e�k�,�7��h}��0y<y��"�sZ5������W���4'q��@e
L7FI���_K�?��H�c��g���cM�cA7�J�(6�[���'[2#��;�x]�M1j;�6pq�jٗ�v�L�P~��3�y�ڡ�#f/��}�p����
f��BA,���dE�9e�6�΄f�WH&Z��D���w!2ߒ��;AQ���O�mt�&�3Ax�����׶��w��6����CP���aGZ�鋧�̅mS��&�?�_�
\!��)w9��ǂ]Vh߹����B�zp��_�%M��X$��,#��ce�OM�AӲ�R�}�OMCr��(�XQ�(�5XVP��!��|F}���؛R@E@����I�9-|�,t�$�,Hd��V��}��+���u�C�/��h��`��9�w+C�7GP쿌�:��+�Fz1ִ'؎�ɦ�á�p(��tε�����6%6[�=�'҅:��c�`hn��Pk��w�T���z�Y��|��ĶW���D�U�w���?&�E׏qس.��e�7c�Ch1Ͼ�f�J��&rb�K'K��򛽎.�.�����Z��'r��{�דQ�o c+2�ƌ3�@���r��5�vyw�	�.�:��i7AqA���l���啲��b����#�@l+"����S����馵�]m������J&�P[R;�`�)Ya3���'u��Ot�z~	>O�Й��������8K�`�\��$;��;e+��������<u��P�M��h#���7W�G�?�vC��8�#Q��E�K��b嬤nȕ5	|�\� yh�O��$<V\�(DW{���q�	B��ruW��{�fUA��Q�P,5�6Q�l�D"2]V���n 7��K��7z�Qn�1�a&�숷鯧ݼ��/ޕ��h�oZ$����U��0P.�ADx7� xЊ3�#�
�����I"�?��g!�`�#PѮ�El#d�b4E�81x�-���LW%��u��#��ӨV,]��nb�M�#�0��[e��Kz��~RO��{+P��g5o�0���+����٦�'L�����y�О�<���@>=���^���H�8<}G���V4;���O���+n?ֆ��^���w���?�Fcgy�y�`�{�d�y #�#�~�o[I�.���R1�K���uٳ
$?�����u+TO%b�jh�b�� v�_"�éM��Z�oD�:���S�e��y���L�j�j��y%&R�