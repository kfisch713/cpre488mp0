XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����݋~��:ӆһ`�K����]3-�+���7(6C�Bhu��<5t+[Ժlje����Z螒�3G��oM(��K�!�$�O���2�MC�j�'.@�ba�*"̧�9�|�[]��=sv�8��4$���i�[�을��la�]�ܭA�f�4�&*'^��+k'�$�p��g%X6x��G6���� |�8���1]��������¶�xȊ\E������B^FX��r����{�KPF�Ix=�X��e�΄�3�{���Z���R��J��O�N�����hj��i�/K>#�E���'���%����i=�m��A��t�ω��7#�5�� �+��t�a����!W��&yr��Ⰼ�`�
l���7j�v�ȣ/ ��`��=<��pI6{p���Mm�R�Hk��Nr��7��:kX���"qӄ,wĤ������{9�L8Ԃ�6��;��H�:��Uԩ( �1��»�\�j��a��Wn�I**�Oq5Ց��̰����\2c�l�L��I��k	s��
�g��,���]�I�e�B6���EN�g ��&��Q��|4��y�vR����~t�-=�����L�");�R�nx� (�16@��Km���v���	�A�2"��&�7wd4�U�jj��l��_�cDm�Ɣ�%>��b��~4~)�au2��[\�9od�0��@w���gz�{Q��t	�	Ƞ܅;�շQzQ�zѣ~�%��Sf�.?m��~$���ʘM��j�KXlxVHYEB    1853     810���	~�c�Zn��%w{��&Ͽg��̠�Z�vQg�d�Y�A�w�[��w?���N0#/��钁��
�O�F+XR>M�I�v�E��J&�|�wv�K)��r	��%���<�YK��@��Q^��)l�ÿ�d�<!�X̟/bP�h�8�#�%O��'�����AJ.o��,�u7L�%߽�����^�!�B.f4��Z�E
�&���\�!s^96ɷ��Я��h���?Ls�#7�-�Y����N��/=B0#G:��&��_��P�1m����9E/�[<�FN�=�M�&��[��+�U�_��WP���0��s�ٻ�Ǩ����qp�$�t�)-�W�K�8$O+d��@k:�Bcէ_�d�~�`��UԴ�G�G��8M3����<�D�X��iWr��K�)�}��we~㺜���tJR�yZ��{�$�v#n+��r׈�W�%�z@"c�uj40���ld�o��m��	�#�� �޼i�+m���=�Jeq�4�����#��aC-�y$N�*�_ @���l���/��]�e�2�i�8 g��]*�1�O���-���ة�{p����Y���VH��ŜP<ǀh2i�X(���د"�l�~ĖHj;5����+�� ����~7�$���W�qd����$��P�����"j���,&�k����*��� �h�G�������hB������u�_
s�4,�����A���a��ё�Y����>/�T��K�VA�V	Nc�hu�����C�����DiXι���ܪ�`�-�hA#\ִe��[d�2�}��0<lfb(����2���ցXb}]���2JҵI��=wU�v��	�z5�(��cD�{p��vv#m\���=f'���X��E��S>P�
�K�v�9*ZAَ�ΘEa�劋qX��^C��d�%�ކ���0X��� ϱ��WA-�� x�s�ps#��'9n�]v�Xzך-*�>@m����&b�����<�2Zq�����Gu�#ݯ�e�]%��tmlvE��2NӔ�I�=�̉��Y~h�\1��ߏë<��zxDĊ9���� �D�����������@.����l��8������\�ڋ��?�����Xꖠo��6h��$]�^������:��M�������H2*����cz���9�.��1> p�P0���v�_d��|��FQMo���+&�A�ʺ~6�e�#}j��.�h�S�cG���+�" Ǜ}�<� �Ӹ�;��aS��:]�}���]S
!t[��XH�7�g����|ݥ�d��b�(�*%v^ �~���*gg�uō,��T�ޡ�A�-�3P	tzi�ΙNJ��=A�-�W$4��a*Ե)&�S�eD1�(T�S�/�P`��Yx�yp�#���+$QrVYF�j���>d�&]��4�oϚ���];��a�u�")>X��%��9� �aĲ�s��"�m�eKf꼏� ��1�*ڙ���y^nm�"1*�>��gv�E>���+���@��.*�i��z�U���u���g��w&*�e�5]�TJ��>5��r�ǈ%�P]ׅ���gS�z��}L�Z�ɏTw�vr�{���}�H���M�$�`�0�Z��
���B��� ��8���^e
�y����1���\�]������?�M"�EI�3�_�H���u���{�x���\�q*i*��6��
H����紭PqV~k��90���6V+tj*��v�d���3�(y����|_���z��7��Rx��P_�����M�LkG������Tg�Q�ϴ�«�-|R&}���6�М�+-�l�Hv���_z���m~�f,6�Π�O�o���Ҷ�	��Y�M]�Ŕ�R�4`�?���m>����<���M���ۗ�l�L+��j\Z�w������D�kc�,���s�Pe-ȝ�;-T�b�Twz-R^M|�.���GIX��E��b�6�""���L���q�s�
�%pjbe5{)Bu��n�B �;�R����H��~�i�9ϴk�A�\�e5E5��?�8
�k"|F�v8̲(