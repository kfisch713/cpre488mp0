XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� ��p����)R�]�+� 6�۟���$�?(�]����7�v~���u2�aD��zݥUf���6}�уSQ<�f�rf��S�i�%��j]�{<��o4���s�P6:�X��s�D)n�HM��鮣<a�V�� ܦ�U@/ߊ��(v��kc��I^�HE�r��A�.��P�5cI��?�^���f�^�#���01c�/���`�ϛ؃Kx��7�W��Y����H�-Ϻ�fb��;t���0�С�B`��W�3T��\좯{�չ��W *$�ߜ��� ��탎�x�t,���:�>+�d�c�Xn�- ���[%cQR+fm�F�\a`��Ng�)�����=|��N/#}əs ������'�����2XϺ}W�����r���y�԰��EWr�pbnB`�c��b'im��S�f��<.��zH�m��Mh��,�8�&{�u Ed�?M�t9��Ź+�6 ��Q��[,}"Ĵ�_WEA�>=`�ӟ�ҡi6K"��čA=F�V=�xeaj�[5��_�U�-#ý�|��43����X�ڈ6i>SjQ��HW���>���0�yt���4lSdzm���W�w޳�w���Z�Γ�(�&gv�&�FX����>S��rt}�Br��3�%�jde�

M����n&�&�La?>�0W��Ej���.j�*ڭ�5s��3W�$��)�$�tb���wť�Ҙ�e��W`�rmv���/D��Bw�d���/Wn5�9XlxVHYEB     f6d     6f0�16^�C\Ib�z�-e�pC�d{\)��S|�
�2�OC>T@FU���-ڜ�AU���0"�;�]�m��"��N�š`�����\�,�2v�J����C�t���\��*>僟�2��������dC�E6,�A��~d�[hBC�t�Zࣉ#9%���hMC��*A�\t=Ҭ�����9�Ś���"����P]��̗��	�1Q?�e����u�{#�%��x��6f4�MG�kb�|e�&�yG��Os�|��w�4B.�`ּf�k扡� ��T6 L����BN�5(ŏoA���:S�-�	pZX��V l&���)4D��<��?+��=�VX\����h�2�_����ո�WvV��"#oz�:�����ۭ�6���!w܆����j
�1�)K�2�����֬HJ�]�k��'q��C�̪�ɡp����E���|F��&��4��`^栌�|�ߙ����Vr�A�\0��~�[�?�!��Y'�x�ONجG��&�z�(Df�}�*z�x�f���h��	��EӢM�]p���{b0�)����UxQ鄦fs�^��I���=���GM���)��0�#�f�<�9��U�0z|�v�Ղ7��̒����q������\�*���iԫ�~K��H�*��=��S}%������y�,�9��������漢�]��~��X�,�����r\�rR�*���D^%����/�w�@wh�P�X��hT�ӫ*:�rT	��݊D6�9$��T����I
�Y���V�?����3B�����0n���t����h�(�$�����3ξ)�'����<5�]��ƺ���A��`�[���Y(�����÷9�e�0Q����b���y�'��(�a����}j��H!2@$��{}�����ja	��sN�1�W����FFn���i>�/��	��D̈2��׮_�&�y *�&8�'�._�]�u����8,�Rd��'�%����ܭ��$!K��9��^�^�{_�<[�7�(A���<x�,��@����yT�{�"��W�Ӣ��T�ֳ���ܩ�w@ֳ�~'����]��z�}l4 �\�cȺ�L���T͠F����g����u��6z�!��K����*�]B��[*Ed,�Y9T$Nb�����Ok��A%L@u�����#��՗Q���wz~t�Qd|���q{`d� a�UDR��<c� ���[/c�>�Jwv���K���:�	in�8
.N�e#0DUr�!y3MZMf+��A(�I�/�vzK�d"/����7��Nd�!��ȭ��][(�Ju-4������_��.�^��UO9�]0�5ێ���kaz��kQ������0>)<:��fO�q/��8�V����4[_m�D����|Ѣ�Pj3���Z|(��'�3Mc~0���¦���T_{��)l���oX8� s��N��*Y=k
�'�dH���+�(��.L�+�\S�*��+�Ou���)Tf�`����C��/3�rO[��Jᥓ1�1�wh�:�=$K\'P6�%I,��<����(��9_��
4��2�5!���v5�΋�`�4��-��4���X�D�$�Zή�K�~�f��e!H��ꡄ�b��$�P-,�+�����B閬�6��<�a�)6a�.���X�}�Eo���+t�u�&����ãRk��.o���� t8z}_��b'�tQ/���)�&O���

,8NR�qNu%kf$7�^�oգ�B5MLi�my�]5�