XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������'"�Ƅo2 �J�܃7�,��ٰ�1���~�+|�[9E��ƴxS�dcaz@�MF��f"�K���L��{k�7��)���Kk���Ҽ���v�
^8�O��P�]�+ 2*�Aѭ]^�����h�c�����)ɋ��^��5�+�;$�YNA��_S�|m\oIӒ��*�Uk?*�ف�>��/���{�7:*�m���'K��Иe��
����2��ge/뙣�#�ċ��ͦ="�3���ϭߠ� j�����/��?����>˼7n!�"%�K�aO��_������-��`����MbĶ��i�B��vow��uˀ�:q(�w3�o�,�Ҳ��6^Ҵ2Ul�7r��@��?k���Zs�W�k6`W!��a�adU��
�=��p���y�^Y�
��>�� �5�Ս�m� ��ND(n�t�wt�mc8/���(�F��R�����@�W�)�O>k/���IBz�d�V�C����X���2����Q(�V���d��\��KC=��S����/��I��u<���W�҃����`Q�M��GN�`�@}�b��D��\� #I�r�^��Ī���Xj�n �����0���(KEu��j��4��d��B��Ǆ,�T:�&e�����h�>s+XN�?"�2�#��Q�h �,;��{����b���'�eh��x��6��U1���+ �����s�x8y����б8�������]�0<K��8��au���V/��a8"vp)6���ՎTXlxVHYEB    b3c6    25b0�$x�&�|x�X�^nLY��X�+��O�gѮ2!�фiKj	E؀�H��C�ǫN�0�̉��>
�e���Ziw1%�*HJ,>(�03,/��| �,��"�a����u|�"�W���������Z�,��iJ��Q��?ܬr{��*����Zn���h�ƺ�iL�G��C�.�H/m�A0�|}F"B��)��n�v&���PD���jeD�0�{$�
G�v�l-��6�A�p�J���������Υ��䜲��������_Uy"�x�"|ߚk��uL�]L� �U��6����*:�.Y�&í��ncx����*���W��(�0�����i�xw{�g���=�ʴ��
7�9��>���Ņva�/�nM���7�4$C킹2�G��&<��h{k� m���C4��I������;�dJFBS:��S�X��5�{���2\�3��=6pxZ�Tk���q7�6�O��pLjg�~0������n|G�A�����`�I<(����79��"�w��Z�����ѱǾ�������4������;�{�y��h�$j�`�G�O�;��` l)��gĝR����`�l����3�x��"�O���ggze��s�TN��/�>��1W�6E߄6�����3�S�d�Z�d�nu4ͧ�M�ĸ^�j�;PA0�7��NY�*3�����'�aGS��P9Vʬ��.$����S[/!���5�-�|���p����:�ݿ������ �3� hg��m�Ch['W�*��[��!7�_��}'�r4����#O �;�]���.����{��ol&��χU�&}=&�M���HZ�E�R�SQ�XMV�db�Ҽ �&H��~J0:�R�?���=B����a:�e�tuS7�Mh���M4�>x�)拞�c{��b3�ջw�J�K���Ъ���|�����S�)/?Hp��4'�����1p�f��TV�Vq����[�k�mx���U�<���W\c��a�yɌ���]?��4�$�ueR�6?4�j0)ȩ���<��Zk�ӊ4�����Ze����
!o+�}�Tu�o������U�oo���շ��9�D��)���2K�����a(��g��AH�;穈/]p��V�j��	?U)=�M$��0���:,Jp�>	9���tkn��-��g��{�Q������}n�1�Yj0��Ī���a Fb�g}�����C�k�BnRw�O�N'$��� h[�m��ī����"�����	��_뜨i�N����/lґ"���"�AG�t��.�"�`�������i)�~���H2��U��(k��Zx:��u��Iӄpʶ����W}��thB�`LN �a�����3�1�Y���{9w&`s��I������,�ݕ�;��%�1��~��̓McΌq$L�����W1��,W�ɜS��"<�u70�5��H#��W~!J����/IX�u�%[C�`�1�S+~�\�-�ɽ)Q-�u�$Ȃ�w��$�  K��P��M[}�BA�a�|8���H��nJ�Y�%�E)�f��#f
f�B$��٦�.�q���v�5_����9���d�i��XG�+�����.��|��^kv��o��obm3��;3�_���\cc@�C"�r33��Rh�c�i��p�T:F�h"��5�E��
MBֶ��p��A��x�4Z��K�:���5��g�����S1���oZoP�{�UE�O^}Ll���3u]�#�76��oƀ��z}qS1󑤤f��Gf0z��q�G�ۢo�\�$���t�ͣ\���D�W��	�Ye�)��VS�.~�b�	���F���f�Z�Y�ث>,ƌhe�����e��X+JO��M;��[\��S�����q�N��Ӣ|3��I�X�����lxS4�9�)��o����x$�p�>�|�k*P�r�q�����6�Q��_�*H��BM��4яً�܊&;k_�3ĖI��KT�4f���=�C�~�*d�jq�V�Y�Z��y�q�6�)����U�3ˠ��a��y�*���+�N�����L2���ȸt�$�	n�W���fG�|�ߪ�o��<Z��x�u�"��;�z��yN�͆8�Q�iY�Z����1(Nl�~�+>�� ����>�Nl��0D9WP�� �W����N��K�E���U�o��X�;j=2-q'�(�������3����m������D�~�E���`��@���nk�F� G�]���ke��N�n"Au>\\Oqu7U�LG�x�mC�`F��1x)�/�7���2)\a��n���<�n�߄����2�/�UlE��������e}��Њ�+_T\��&�r��H� Z e�+�.�X�)������(U6E� ��P��@E�!t�1����J�J���B"���KM�H�(mS���`/�
 ]u��̝�t�\�K"r��<�esc�z�Y����a���_F�>��7��f8��]���ed��D�;�,����CO��"��~���?A��i]0S��!#�]��	Ƅ%�P3b��i�z�ܕ̂G��*���7�Kx$�1o��
�%reH��
����w|�I6(B�����?�^ji��PS��=�����q
ֶϜ'%����"^1����cU�P�e!�5���=�	ڻ܏�9 |���Fp)l2h��W�{���۲���$%J����WB�cO�Nd�U=����g�g��7�^�Mr� �s/� ���Lg�!�	q��f� V����mQz�
�pv��s{5�Vjy�YZ�5-"T?�������ަs�Tl�
��+�a�~������C_��(#�W?�	��)�,��72h9Vȝ�b���+%F:Y1��$��n�B.}t7*	������)Aa�[��O�(��}Z+��(�K�T0�"�:��M.�1x��OwPn<��k�Q�8�3V���i{F><�KD�����a���#��?��������]ј�n�)���d]E.��a�x��� pU�,��bm���o����.��l$]�no�Ndh�x�@�	�`�5�v���+�!��:we���&-�gG��	���z�ûm�טΎ��!&��(9�m|�A���t{��ғ��
��̈́�	g�7Y�b�>�BO�v��{��� �QyL�g�C��m-.��uY��W�E�(�݄�WfRp�z*��ʩ4=�w+Bzxfش(�C%��ȿ((�/j�J�i	���x�C�Fk��5��ّ;\�zJ.#7���j۳�c/e�w"�a��3�XK���A�e�������sq�"��b�|L���!'�*H� �<�2��m��=@�K �O���5>b��_n��
(%�.����'�{�?�2�7&�����0w���������Te�I~/^�n�Vh7d�QD�p�Sw��!��2/�B�V���Vv5�ﴨ�;z'�f`��i:h����� �ʾ4!�Za ��X����`\���:�Y�jڎ�=����oM��ͨԌ�=\,h��M_�fJ�j|�D��4s�[�jeV+%6"x�Z����{l������3XF�!C��״5p��o���H����":CL0�K&#`�QQ+�`�3��/��S����r���)�`.��U�$}�h��*j�Z.
PV1ɕ��oS�/i�NV�S)CT)4�jL������M�}~�a<��5S��o�7���=X��_H���sC!����-H'��"l�4B.;�@����0�*=�'(�$Z�P["]K���h�{b�l�p��9C>�ܔ�ؤf�\�V����ވ��8�6�kE4�\�$oJ��;s�<1k#^���gy.�]�'���.��V�v�XZ�	{�k7g�,��B��`�n���[L�Ei��f�������yX���~R/a�%��kZ�U�	��]��e�^ʰa�_��Fl�S᧥��iT,.�"&,�)�&�Y,>ε�ىZF��Yh~'W���{���uwuz��( k�
��Ѭj��D�,�䨤n.��E\{6����Am>�������?�}� HL�P=@�9�S<�0��̗n�X�0!r�8hE�z��`��I< ��,���/ ?�o�8mp61��
_̛�7�?]����1Ag�-}�;my�!�Qy�|�Ǳ�ӶI��j�l"T7��&OPn�{Z�F�R&���Ӱi|�>X��;xZl��3�����2��\g�FWt��R7�{�&k�_g��?��[�:�P�,4�D�9Y��v_ņ�sird�T\ǜ��,�"|䲾��{5��ϝ�Q��U
��D"�q����^��g�"�"r��[Vm	�)����蘹9bj����:A�־���V�nvȔ�� �.2+"Ê�e�b�Ô����������S���W����r�ƽ��w�������]a��|��t=�ѫ��P>'6N�! S#���w�m�p+gV�7VĽ"E��C��R�3%=�2`�̫(���y��4(���e壂%_p�.,;$�[�%�:cBZ�q�p���z$�|��&Ď:�)���{9�~��،����``��,�r'݇�ː<Դ�P�9�N ���y�8~\�ʲ�+��q��`��4;���%��䢭���z�w�X�ZZb���)�S��~S�3��g?d�<0�I��fP�jX�[�ɡ�Vu'�8��1�F���IU:C�D�qް 9:���~V��|"mD�ꪴ��a�C�L)�O����A{�@?9.^��|�}d���Q�)�A�B����k!n}�i����W�����wG��Ob���=�/�1b�7���,,0��n�`I���@��u�)���pO��g��� �9Q/Z�#�o��t���g��e䨹=��7Nڇ�4�,R*ա��hbRZ,{�U�l�&[۝��D%fh�'��T���M �(��2H�P�����'T��$��e1�|s�0*G�g#;9���m�K'mPP����|7��a��m��=He?2F���sB�B^xip�8�9�=��m�
,��|(���%��fe{�&
3QZ3��S�Ƶ�rhǏ��y�'����Iŧ0�߲}��X~$H��jU�y�Jr���^�\.5f���lF;�<�ǂK^�m~Mc���ULBj�J���SZ���k�s<��iCƱ���S,��Y������'=^�H�VjҎ�����^C�W�aX�/!���D�,I�86����t�i�Ǟ�ۍ�)�����N���e�B|�A6j��Z�
@���y	�
�0ԫy���Um�e�Bmg;�E��F�!�n#��7?Y�b��Z��Lq%�C:�G�-�쫳����j`>��v�u=2P$�������<2֥����w�1	c�Q\��.lO�Zj.mM\Y���y�t��\��}�`����̈ ���SV�$~m�K$���u�eh~7�&���{�@z��|�"����?�($���]:D!�?^�C��]��qiW���6+��Qhż�vn	g;Ll���[��SLB����#r �������\bѨ�dR��:v.{�;lְ+��}����C����գH�p���j��>�g3u�`J�Ͻ9�W]�G5�n#T
!,1��h�%^آ�v �W�����tYG�ݢy�a Z2�����O�fD!�XW�"�08-���胇�GS���x��?��0���C�yD�u��Hj*U��0N�Gu��o�O��:��6U�ҧGX]B߳5�fH9͘
$��[Һ��8���d�y7(�/�T�����2lՊ:O�q��\��8��������G8Ͼ��-�$V���ϯߏ��Z�'�'�-�e�0���sH�7ǐ�"n#�Nͣg�Q4��ܸ9W��,O���i�@��ڗ�_��Jf^�d���8-o�D8��oԙ����I`����&*ߵ�"��?�1m�l	9��3��캾z���/$3� ������V�嬡�$8bH��W��]�E�C�G�!M�yt�6����ӧ;�����0.I����-}d��-��ɣ��ݵ+k�I���!枓�������3�'�)J�L�ö���Ȍ��B�K{�s��K
��n�#G��[}˿Rl���J҄ݏqT������7U��u������+�zX�4���:���c����H�II/�?��zH��x�.3�����:���ɂb�\$�l7
�{t�Y�N��#�	H w�g�)��|?IP�w�@qc�	S�b@��#<��h�6A�m���[QL����〵���=T "X~Shcސ� ]\v�gR�qӻ,4����*qT�#),����pzC~�5���$�6��Q��~G��?k@s��+F�F�,m��������þ�>7XJ�5a�oOD�{�ګoU��d���р�}�����"]�i6�9#f�8%��'�=���.D6�@(�ᠦ֧��� ��l�1���$8��" V��C��Sz�J����
��h&C��T��Cc�g%Iɣ'W
��A^hO�^,�,*a�^գ�?�1St�S���N��R�
:�R1�eC�B�=�U��W4k�y�xeߦ���m#� ��w�EPټ�kh��=��l�>QRW��@���/I\�M;�#e��h�
`U��p��	.�����M��a+i_į�߻=j�थ��PK֣���S
x���|O��G�R�MJ��]�b�%�`&r��Ŷt�zy��۽�,C5l&�W�*�ю����sB%��
#�<L���P��<�*zY}���V�ו�I[�#E�.|v$^Hf�8���=$���v��_��3ر(�'U���Fs���������s�%bD@is��Lfx`�8 j7�$�u�Hw�������B�b��å;���&��➭�ңoЦ��+b,ś��FaY�-��q�͋��w���笑�b��7��mC9�.�z7�!�:K�6;�[jm���o7%G�s����0��m��}��U�U�
� c��վU0��r�m�?)�kG�K�p���5���B�Ե�vI.�����5~�1�:T�ccWԥ����~����)�@�=�eE�1� W/F�-y<n�HK��lv�}��se���nRLj�!@ߴ��-q�.�o� ��̦(N+=���7�.$�?��!s=ހT#�ǘ�b#�����h�KB
e��l˝`�!��.�����0�5��+F9)""����1Ѳ�0@������3���lo��q\S,�A�2%�ާ�)�Ц��.0�}���#+� G����7Z&	+	�Z�~v�=�.y�����=�.))��-F^
��.DRaf2"��i�lp?��(M�̮���'�t �W��c�)���N,]���h"�������e��%&2Fd�w �����j�d���{�ٺ�.{�V�e'����/k
��[�6Py�v��!!�[�:�`���E�]���c�$�ˤ���x���]��{�W�x�
Ɏ�q�iw��:[��G��5wU�>`�ۀ����p�q����z`�C��Ad?��~�@SF�=�Tˑ��Y����D���dpW�ϠFhñ�FN��oę������K�N��x�E�����۞q��h/I��We�Ӆ�f��*��ҲѥL��f�3���r��3"2�t�ҭ^�ٞ{��#�[�j�0�,Ht���u�)���؛�#�Â|�U�(-y�L����q���73˄hdS�z�Û��ς���)������q�|�#Q\�qR3J�4��X�0���xt\��&rD�F�f��@���4�xv��1����� 'M�y�?9K�����p|K��NߴW3�}^Q��,H��B
�k�7���^�׬ v�R���xS��\f���Q1�0�͖/Q_���zBQ��Y�����Bܸ� ���k���hF��&�����S�P����ji>ЦJ�,x�UxǙ���YY���K_�J󮇇_R���>��q�p �>T~G��c��������6p���jzY���_�������� A=!o�c_<��4���8:c�hL���3,��N��5��c�z����TG�9Zg6�F�����1�b&�3 ���WM4C�C}!hh�g�M5"ʌ{y�¶U,�0��ؠ�
{q��
}��2���0Ɗy�Vj���PnB3��w���x)4Nn�N5��~����/��>�m��Z������j�yoIa=�AN(��{{��iK�W��U����B{@N߆�\^ t�\y�k�yCo�� o�t8�,�[1�d/�)�����k/�.�4�N��E�/6�8{�Ȱp�"&����# ��/I�^9v��/-q�˝�(�L̫���L�	ّ��蕬�@��]0��ܑ]7��:>��/RZ[����ԁ�� �0�)�5�[�G~܆J�)���$�\�v��;#Lۇ�����}���伲?��Qd%J&��^���>�Rxr�Ӟɨ���|U��E 2�%(/�m��C���#K�g ��'��xS2GJ�2}��Yi�)�5_�1c:�����q"9E���J���ڃ�:I�`m*��V���LRI���ıڒ�Q�W��ds�m�Ez	 �����g9�a��jR�o�[幆e	V6xK
�+1��2���M�#O�R0
�||.&�+,�ؔ][__�p��m�v�����-�� �;�iU�����5�}@bg�����V/��!�Oy�B_�Q-�a�d�j��[ t2TT�& X[<8�����G\�H�O����P��Tuҙ�y��s�9�4B�Us��^K��n� �>c!��(�.����Ƴ2��H[l~Û�A��	0��j�Ȧ?��ۘ�7�rb�ޠ%N�T,�����:Y?#��5�^>��Z�k��-JŢіE%2���3��3�ф�b�1$��I�K7�9 %�+��^��R�xd�~�%g�Rb�^���x����W�����H.��d	�)3�&)�u����ڝ�o�t����j�p���Jש?�\׷6R���2�oԧ?p5㣶1B�e�7�U��L���")`U�jl��{9��9����:q�_	ydù&�#gHU߳>2F)Oh�˛Mȓ ��wpҹH��gL�%�]8c���5�����ϾG����$G�&TO/z�/�=�虱4;0?/��D����'u�V��b~��X��Ԑ���O�7�����E�w���8�0~�N'���@h�f*}8�r~�^ė�_�jt������JV݅JY�)E6�z�Ort�/j|RN�~�q���菌}��p�7�!��F�� ��m�.�	��v^�v��D��m���Ԗ?�W����u�T�qaX�3�ܔ^���Åi�,��$ki�aCɼ�n��;�Hq`[%���nN��}stƃl�Y����`���a�ڔ�0�w�x�+���tB��5��o�(�5�,4��L��y���]������~Ɗ�n�-ҋ�VU���S ���