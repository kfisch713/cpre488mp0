XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������>�����rBb�9퓎���m�E���]>-Q�CY8���$V����UF �
1���Lp�R6iX�`s)���Ds��4D���ݵ5���Q��6��l��o�����'��wro�aLlF�fV��R-�n��0u���gu�ž���a�t��U�#x��f����u�r3�Ǟ{��B�G|\T�������)�Ѽ���L�OFޛukd˵��й)r ��$�3��1�P_	��ʨ�ׇ�U�;e\K��n>���v��ݻ�"�$K���������M��4S:���{�]8����-^�U8���=	��S�mi=�8�e��h�-��I{ES[�����L����YKzd�E��SU ym-s��2�_�i��xY�p����!��W���)��U׮`W���i#.E+��,,ؾm=�I��ko�'Bj�`�%��㐦�,�p@��m圿	�5r���p�йQX��+�|~rZ>�{��c4�ɸ�LR��@��ѓ�Xۄ�{�����!_�5
�ff�B{g�&D��V��Ca��x�z�Sϡ���I�D���֙�6
�"jSRf��r�1�	H��Z�K���Y��B0wԃ�g`e��FΤg���%Bv�(�#�(9�� ǀjHק�,1G���t��n�V��Ulc�Le�%�5ӝx'B<�E�ۿ�C,�1w���n�"�t󦐦��&�SQ�K.��:o���̭��^ԧ��sKu��\|�:�a1����с�f� ����/�|2/M��/QnXlxVHYEB    42ae    1110����5^��:�Χ3;�O8��������R�����袔�M�1Ώ�U��di��/ʍ�������uŹ��v�U�)������l)T݆~��dg&:N��\�!��&��-� w]���#��{0>ۇ��Ӡ]��<��{��+^"�/\>Jش� �6�C��w�d��^���O&x)��@T��J�m������]�u�M(ڃ���>v ����(߸/��tLh��<(Ҏ|ȑ�lx���4���dv dŷzd�ȭrJ�2D�G�r��(`�[z����:ze�̥Lcg��*�:�����f��d >3�+�*�*&\�W;iφě�Xu<=P�ED.�~ıuǻe��F�m��*��F��[z0-[��"�x)C���[J���#ɓoK
��v���
W���P�헦�`��I���'t�as���2u턙"f�ѫw�ڶ��=�ρ��B�u�u�'������Uf������!97�/� ��ҼԎ<a@( :��W��!���'����I��d�[ö����ܦ�g��=<��Vk�?]�i��]e������li3"����O��T:�eW�h%�W���֏9�~�7��t�1E�#���"5o��*�'J��5(.\��뼾�V �Ŗ���E�(���� ԑt�+��L����	Qg	��8�7$�
 ��:������<?�7��,��>�i]h^Ǒ�¼S��6�jP���
M��5�.'+��V�C����p�FFI��#�YĄW̟�Mُre���T6�`�!yj 3w��؊@�o�8�&�%t;�q1���߉�C����#L�u����'T�?|������>��!� ��x���!W�,��0=�niN�v������C�>ȧf���?��1{��&�9|�+�
щ2-|�"�#y����3��/��TϪG��ԩ'3֕$v+����:�<�,���>�Z��]��gU6�R�l͝�:������4� �b'����,��;�b��wJ:Ӂ�rY����|�rY���F���C#��s��{yO�+c���C� �РB����Ť�\$��&`>�=ǉGv\h.�Y�ke��W���?�T�5��E[�tq����u#&��,;�~���s$�Z�����/od�����24�j�����G�	�9�'F�~�������.�IfވܿL���Yx�.j��j.}6�S��l�f�9��U��@�ߜ)~��fP��#tJ��.0z�=�s�Շ]i�� DNc�w��br�2���@}r�V�
����_#H��D�;6�?�@���Z���<O�?�$�����ȯI9 �ώM�v�Lv�������y14��;7�eŖ�c�6��ŶQ��7 �~V.r
u/?�?�L�k��\}~��BK�\��m�[B���t��"���	��NP��_�^5D�f��q,DV���5�*Xm0m�I�T��~�~��b��F�'Joo��?Z3e�%�,42�ЃB��s����s��� V,��.'�������*�*�}uM��tJ���!�ܕf0L��#5��˲��C�mR������_���B�d��)�Y��Z*���~��|� ����>��ܾV�I��Y��%��S��Vkd|��C@���	�(���a Y|�Mm�pLK�֫k�+����ѫk�I��G\�"n3����Q�"h��ܬi�n�}�ѩ��|��C�˪�S ��E�bFp��Xzk��In�w�f�s��eH�Ŵ�lE�b��2����"��?�������"Jϥ��6��������Nq�,�Z��)�*��j[��2��&x} ��O)�]4=�Ah������Ɓ��CqQ�UU7lɬp3��wA7̡�|�>�iq�~��)R�g0W��n�Y|K�\t���=Q�;����[�$욡s<�����1w9���f??)�L�X�h�2d���3	t��@��^��0�+/��P�5*��D���7ٛs�C&
���)��ǒx��w��W�kN�v�_���Ef��t p��G�b��$�	l��E3b@Jm���;��<dx��8���p���]��ip��z��lª���j����w�s�'���p�����*��o!1�̄�	��{�Wި�����X��[.���P�<44r���ZR�	�&��W�%!G�A%{����~�r��5�@#i|�%��H��Q��Z;�T��ֈ]e��a[�\J���COX�%�@��i��x��ή`v��-b>U�}�\32�s���/�:u�R[��4r�����iZ���y{� �E�:½����(z=z�xE�Oi�h�&k/��W;���NG~����2r���e��k�M�@���('#�W�XY�I~.���)
L���wcKƉT-�P�g��k�l���O�Ԝ�W(���t�-1ƿ\�QCpi�IƞV�Vl�"��b�(�B3&��Ʒ���J��J�r'�x6@tAײ�4�ᣱ�cv����r߷��"�{���,[�8��/����1��.s-�5�*��f�t�H=�H��
�A���J�-���4�h�`¨vPQDhN;����vk'��B�e����߰3U3��X2{|r�
[:�金��ۺ۴~�j�B�x�o���D�x��eNH�!��=�v�gs���5/[��R��ޡe��@B�dYGu�ʱ:��ۯ(V��>H>��h:E_F���s�<�-�8�*G�< �wB?����S��-��mD������4������A��b��I���C�d5�--0ړ���ՠ�Vj	v��,�d�3�]lU����K����Hf��aFGc�E��I�,%�.�-e0��~L�yt�7���I�M$��o0!~W��p��_��}�$0Gy@K�5��9�=�
R+ō����_3�)D��g���5#��.%G������Y��*��ؼ���t��P=A�z�sǿ;~ �ms���1t�k������K�)Z9��mxV6a�Q�mK�Sy��83�$µ�~Ņ�\E�E��U'{��o4�c\�S3dn`��	��k2�آ����׌�:}x�Ɵ�#g���{/�!f__� gH?S]��6b6���h�d�(v۞;�F��ɼ��ՓC�.��<o����C�!�m�)�	�~��3z��o��n������F�J���D��+�r �#�^&v1iG�[��G�9tٵ�WsE_�z��&oO�x{�'#<�t`��m�_o&��N0�u��(±����%h5$��㦽��Z�	<X��e�b,���F�o�rDs�
;�6�L����n������5��:9.���_���{�N�� H��Xu�%zT�ݘ�V���
j��wJ�{�D`��X�!3�T5
Oe���g��e���mNp諔汽J�k;�Fo^��|�6$ ��0��d pT�%��s�3v�Yt�r����|��ƕ� ��}2Ò��c���h�W�ޟ�t崽AT��y��_�ǍZKn��F.rZ��k��p������i5��՜���m���>���z�������A�eͿ,������KFg*��;��w������pΥ@�۳�G$����Z�h;J��n�{(�ΓN4"�w�� ��������$�Ǥ�)��eiS��?� �sC��=�U�nzv]Ur����m�3����#�����l+;��*_��4P�G#&G� ��{�(�4#��w,� o"��Qf"K����Y3B$Cc���
���m�e�'���_�Ciz��Ŏ'��f�ɉd-��h�D�a1��r��T�Mj�皞�'��t�����3�K��G��ԥ�84��}J�Bl
p�]jO'�,x�=>�vAA��'7sE�����G�z�܇~��x�'�!����1�#���b8�:�x݆y��7�~���L�'���$1���Bg�QcW#&9�d{�]p� ۫#�R)�ReF�~��;�d�3Âݛ26��I,q$tʪ�I�|�������AHơ��}:�sV�^��WiNG+P�d�P���YM&\�d2�!ę�13x�N3B�h�y;�_�#����rW}]Γ�	���TI F >N�M�a�yu��S:�� M�vǹ=LBf�MU���w���?�X �~�r�x���luѪ�H�W�
;f}�$'���!g#K������)$��\��h��Ê��yUǒ���s�x��zӕB�4=�kq$�ڃ�v�{+\n�ob��{c�u[�
�3S7���R89֭���^��cg�ڻ�D	rPC�D�jiZfw�)'��R5���y�@�^��:$`t6 ��|#W�E<�.���t�!��f���B3�hE�[�!8L�_�+��&��w���\