XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��|�IVo`�H�kWr*��u��y�o�F�Xr�1��C� � �l(�?A!��8lJCIen�M�kǅ@Np�%Y�>�y�J%<�:q�����=<�EX���{�q�"�kj�u�%'��R��X��}�1��[�:Y�|�cоO�[�8���7wo�$�G��77��}ޯ��,o��BTpA���k�2ֽ��vHt��7Q4/�q�8�����|�5�n��i��9�k���J�\F"|��@Z��Ŕ�5M@'7R��qՂ4��8Cy�h}o�\V6װ�X�D
�/{�k�H0�%M_�!Tѕv.!`�ܔ%^5!�g�*�"<�����e[_�{��o!P 8$��b�4�#����$�on蠝�ǥԫ6t�>��؛�n�ԐD#}�|)a\�;����(�?$��X��eU���F���P�:���#L��Y�3���~,�`�
��?P�Rٿ����"*��	��,��n؍ѽ� ]��'� �<	�E.�����N�-$m�0��T24�׳��r�o2ù^��G���h���N�� z��]���'���R��X!�$ޑ�5 .�Y��ӏ<��AD~3$(�R yXQN���Qt�T@�~�Z����k9��K���{��x���V؜�XO(lx���;�j"b�o]�=:�>#�+��.X�b>�x��V��I"��E/�$��wl�����?��Gg�Y��9b.|&��R3W|o7�bLț�e˜�{1ە?A�'���=����9��gvxW�� �s�8XlxVHYEB    fa00    2040rn������0�H�S�l�}��Ӥ�F*8*��Y��55 ,T�fR@�뷝����W$��z�}Ƥ���`�{j�#����m];|JGLx[�\$�ʹ*V9>oZ07�.��Ή�T��8(/w����3,�Av|�P����UXi���
����e4��L�r���!U���-�%
�Bc�������S�ǥ��kɺ����LZ�C��Zr�pK�*߹s�M��ިxg�t,o��ߗ,9�ƒ��
0zN��GB�@��D��O�7<�-�w1Hl��rR|`H�����첉���4�S7����F`��3�l_$ϑ�K-y)� �(�d��bx��\;��+��J
<L��d��ϕn���.�b�E�YŪ�\ )4���eCB2T��ry:��U����F{�|^�^E�A๩=n���}H#���pᎵ�$��{�6�W;���&��[��eѯ������ %e�٨�Ǜ �!�K_]Ǽ�"���c2�Gh��iݻ��'��h `R����d(�3��Y�&`m�k��ۛ�c��$��i �!�
�%�`8k��Z	[�����P�rG��9�s~����Ӌ_��[ԙUfRΉZʠ�yC�F�XT%�S��"��YN/ ��D�,�Y�� ��8~�?�����aP���K��6}8�
��g��ҚѐQ����<#v2��;/E�^��r��k�.y�tO��M#���ÅO�3��/J�
�#��i1�>�/ѡ6=�"�^�l�.�/P'�{}�:^]يP���q�����59t���.PIKa�`���:�(��͕�u(L99DT�V�U��>��C1�n������qh
��}�|�ڪ�X����\
²����ٓ��.B�n,I��	��<��:΁����($��"}f�(kG�X��F�~�̐��
�53���$��-��C 乬_����6!��z�úD���A�4�����(Wƌ�+@�����*I:�)�b!�TL�iL�]��=��O�H �k���4�P�#�B�=	��ݺf�Oj�郢d��'l5z�0�2P��Ƶ@~ ��v�:+x��v8�.�Xw/kdjiS��)���G��0��GH��jS.e�D�#q!�ȇ��
��A��~}O�6��Xӗ�^�>�J]H��̗�W�Q(� BP�zD1(R�Ɠ�@Q�����I����������u�ܒ;��$�Ć���=!Y@Ğ�ޫ�o����'�]:��,~^�ި�܍F�1���#Rebi#�ȣF���S��&ӽ���u�󭍷���`E?�I
W;��E�f�j8H�2\�?x8>����RŖ� m�h��v���R�;�����p���m(��i��v�}�JX�k�C�x�;W�K��Y4B2.��XV�<i�EO�LZe���7��Ŝ�L�\^��xk��42,�|U^��h;�2�j�4{W��yiГ޷�����n�)c�n����9�>�g^s�sF�^c�)�+�]:+�{�N�ǝ~�!Ju�ą�eNYU��Q�H��E�Dw���*����u�៴mE��6�\g�"<h���צW��� ����RKD�Vr,�CpR���tHz��%M�΄�N�a��Cbmf@.^bC����^�c�w��_"�U�l�Xok�ʼ2���˘�G�͠������Y�aT��+t�P<_GѳqL�y�6o����<mL����p7
�o�(iy:=��+S�mC:�ⴃ{q
c|z0�`��b��t2�z�vrVšLoȏAe4�!Sk� ǫc΁>jPgkn���uKt�`�s��*\o�T\?��m�S��C�6��M��L�Cs٪�QV){�#^
��R�z&L���BI��f2�sDh��ѳ��޴�?����h9����.��TbY���� ��I%}��"[���%�J�94t'�C����I��D{k�����n))�PR��B�fȶ������Ple�v(倠������{Y�Ih:Uv���8@! �RY�m��t-Յ �%���mb�xo�	˙�ύ�X��Ƈ��O���d���Q�$�e�M��dF|�Kև����3~�T "���:wj��o������ϙʖ�&���������ग���``7b��Ŀ�ā[��/@0�������/�}(�S����>��҆�w%Yj��뀍�W΁�zB��f��wo��v��2�%%�R�2Rt��D l���a���q���Jq��� �J�)��RC�q��5)D���=y]�L�n_n1��.;JI�IH~t�����Q�v�5E溍�&�s[��| ���oe[9xtG�Uethh�I��X��N�D|�(i�6��u���ZH� ��n�bщt���S=ڟ�J��@~��k����8{�H"�$N�%�xљ��P$!�_C�Y(�B&��!��N��B{9��$�sT�B���9Vq4U9:+V�3=�{�ǇRSd��P6*m$[�{Vkó�?�^uf�	���ُ�?�M�D���B�yiYx  pU���N�}�)�������P9�ǌr�7��O	v�4uy����4+�Y�H�~�+���o�����Vhć�O���s�
�Wf�[�k����s��,����.1�T�c0�ۓ
k��xu�*��C|��(6�������v���V9��EA1- �f�u�'�3>�C����a�<�?�����ڌؓ��Y��G��z�����Yc�)���N��6�/Aųj�E�ʑ�^�srR��CHfc-S-)KS�E�R���'��FZ�z�t�	e��O$��2����2��3���C�JN9H����J��7��$�N��w[H��O�>JC\�Y���9�M'E'�g�n�V�:�΃�W"�4���W�j�iHW%[_�Iբ<y�Uh���Ob��������u0�FO{�����Q�#αP� hC�쬝y�\���G��$YPG�"��B��cf>�&��V��g5�b��$�b�5�n���;g��P���'[�nq��f��x=�m��x����P8b���\����*�0f)·S�������M���5]"n>�Q��6C5-��N�Z�\\߫�e�J&��0��~�w>s�]*��{
�ѝ����Qi�h]���1#d�q�cX�_�{�w^}�:���Z�'�\�/X�Y�lX�s�B䀫�c��;��<3�^y7�Ύ�h���^�ʖ��MyWaJN���+W��YL�sa��
w���"x>
�W�b�]7����{�����XҼX�<%��7�}`�ٰYR�O�*1��z>u�@V��}`����!jz�_2N39�V2�y������C��h���9ȷΥN ���Z���C�*��l���.A�g�
���[�/2&��%%ܮfv�
���W��2��~
"� BqKq�H\`@G����~��ջ�|JU�����x~Q�Sˠ
�� :(X��$�G�'�G_���ni6��5U�Q������9��(�)�ǽ����gRSɜ�ܦ�B];	��e���j��ʥ��<)�{Nx?��QHza�PJ�x7!��T�zM!�y/4������&n ��tl�~J��p����w� ���y��Z��h���$P��aV'hK���K�0ǐm�DwL����4����tZ����s��J�Z��6�6c���UU����k^{�|q���#*;�c�;�����|q�]����Z8�TU�G7ǩ��7a�B�R��F��6��<�f��-}Ԙ�s�����%���/R���+���T87{j��R��֍��9�u��B{1$�	��&_��9�&�l .6x�%2��Qи��҅'�5�m���s�i^�_��S��"a>G�Hm+��^$p��[��E��؏���$�1մ6j�{��4{�п�������@���n�wu&�x�m���6,$��m]`q�&�Qߔ�d�V�o�#�r���/�բk=�mYO/ڗ��&�n,;��ڏ`�5t���� �<VI}��h���sf�u
B�f�>{�6�]o�{�HDF�U�O�=诿���������(��,)�B����/�̗�J��fX�N�6hb�P:�|�XAi�܁����U9Ou�춖���&]I�)����}�mh�h ��ݡKr!����B~�� LzФT���q�<��G;�t�\�2�+����:�*���e)��w�NS/L�ۏ�����wuR�Ӽ]�f��!@orv$��n#iA/LBM-�s,��ٞY��R_a�D�[�TK�c����s"o��E=�}&[#)���������E����H���ٱj��,�\������ؑ_]�x��ˠD<Һ��g��1��^E��|�9����r����ϼ��RW�K۝	�紷�y��fZE� c��c�����r'@q��K/�u2�^]�&�!���2Y� 2�Q n���}1E�\8�dhЦ�̪.���r���|�6��"�Ź$�R��A��#�)�~1��M!^���\��z��g&5�R�&�h���Q��{�w)M�G���i��ܲ�+0�w�wB�,�[� s�5#��[mX��Aɩ�[�ߪI $���h�e���U����9��ܵ��TY|51��P�Р����v���h�.]�?!B�q����\�\�VY�ʭi����4 1?;d�Ջⵍ+������*p؇����K)r�]���4�?q$��t�8Q4�����<�o��#Mc�'�C5��
�G�?��-�d?��M��YߐU���VC�����3�C}��{�6IXY����ےL3l�*e���2�ecG射)��MH��%���A���\�%�ggKfu�k"�QP7��F-9��W����5�TJ�L����ң�}i��Cr:��yh��掠������E��d�m���HVw�W{`�3�� {�p�����I��FrIu�9�6"(� y�޶+�2��QG���!��%�E�fBt�^'}a��0��3�>�!����⿏ya��P1��8��������}L�7���;�-�^aОd�@X�fEȺ�3rO��G�}v[S#�`*0ߧ�̚T�8\
�j�i�! 	�n�R��/[����{��S�8��Ӏ��#\u�8��5T|��
!&��k��ZG�Tu�0>ej5 9V2e0JW�Au����z�h�ĩ���^KER5*��|ev�&v{D��x�m�Gi�kq�X�ԩ?�'z�]��<ѡ�ü�zo!�^��ޭ����������m����H��=���m�*�]d�s�YUh�nFv��+cJ�D/��xI�񷨪��e�*R�~��/3D���X8�y!v��b>�������>8��-�S��Ue� ć<,�Ͼj0�-�GŰ�ڑ��_GY��*�[PYU�s�Q���ʞ��ټS/}rF�(p`��R�E��+��y�}�����6ɱ���F��Ӛ�����wAFk�da���E���,֞Ł@�ۢ�*@�����1�ǣm#S��<D�%�	�f#sz� �b���y�%���dF���+3�ɥ�7K�?��;�	����@��Fb��Fы-~ժyqy&ȄЃ��	b?�g\'�`��)�O�s�:Kװ�	��Ng�_���Mk�h�6|:�`r�,�^+�q���=��+�ui�kT2e��~Q&Ӹ�L4��ǿ��Y5K��i
�s��K��:�p-����*�����Λe�����&]�`���׋�yI��6��dB����qwD�_Q�#�:�΄�`6�ꑌy���Նj�I{h��⼣��i]Ы+)&�N���*�F�6��v�1�����I9��]E���UZ��!��6�B gc���Է����Ŗ�L����:v6I���;tu�9��}1e�0�y�>3�H���qx3Fk�Hgku�Q(_����.��0a��
k��ъ$��Ž�/��Jj���*^�7���G�f���]y��ذ��ྊ*g�&� F�K�f]�WDc׫��d�,Y2i�{��5Q@�
0�o<����<c,l*g��;�r=E�2d� ���+��#w@$�x_<9�瀱�o8�2W��H%����I�� xd�*!�#

��~\U�����X�E�fI��в��Iwf�� =)�4�M4�W�����x�~<��5O�\��STC��XF��	Ģ�)��\���!����Z����Zή.����j~�7��������?��n^*�h���u���Q��]�����c�p�/F��2�y��Ug}�"��D(�w�a֎_��?w~v�k\��C�	<Uy���+��O���G�_�(���$�]M_|���ɤ	���@�╱���l�&?.�α`����~�w�0�^��kHԣ5gz�yt��D���:Vd�Q�>�TCt�l��㈪~�;o��P5a(��f�9�%�)�M�q*�p��&R��,w�ia���d�ž�fp�7�/�}$B{D����^�lT7�n���񇜌�"i����r�2�h��I 3���m�ݚ9%�����4��;W�Pm��0��:��s��0�}h�ߍ������(�
�|�'���`D�y���,O��[�(:&_�M4��Z�_΃Η���^��������e�XZ�g�.�(?�U�G*���eR�Xd�I�1�ީ�P4q���>voU<����VQ&׊���%�uA�9gؾ�� ��+�ڰG���C�BЁ<tƊ����ct@�����b5v�9�U��+�~{a�H F�q*�T��9�A[�Zҝ�m�ٓp��g�/���+�J�%9/�`��T����m��v���F�v�1_���b�\O\O����l�������	Z[���>��Gtx ������!�um=U��*��*�{���b�7r�6���d!*��?�d)��L�P���.���V$��S�	gK��"R��=�]^bH�;Z7�+�x'R���I�8�[pM;ڽKB�
�bc�%q��>��kf�\M1�%9�<�zR���������	}V�gb�`b|�ID`�B���N[�620�AQ���R�%/,�>��͏6_k�/��L��������o�H��{�9��oi���.����P���!��bH�E�A�aT3%�VXJIG�2�mb w�	 XR�i��ֺ�C^Al\�Va���/�S(��ڣۣV6�;�M�/@��>A1|�#�3��00x���Wn�(�w��Hl�j<	�V��I��t���03��0=�9x�z%��t��"�!�U�<��4n�_/ѶX��(M�3�[�)��(�3)fYN�a���7h�	4��tg	0yZ� $�bc�?`��:e�E�)������C����Ա�n���Gv��~���k�-��d�1�p![�4��'��69�T����F+� �Ou�Ӳ.������M�G��gzbE�U0�|}#�&1�bAi���!�نV	��z��ŏ{d�!^��#�h	c&Y!�t~��2�a).=4S��(H��O-)���qߢ��nP�=���9���k��'�
���CQ��t?��;�U���Vu��=�YJ�#����;~�����8sшL�0M�5�
rQ#�$=�wmc;�.��y���k3�tKƩ�5�n�g,���+���#C�U �X\L��.n�%������'7g'�>C�v��"q��)-�0��=jQdq�KO��U�q��9��Q�y����z����r'�߾�$�s������1]�K�47Afj ��S��\I.F��?��FJ(^mk�3N*�,�%�ϲ�h�jXR��Ou0
ᗉdI9R�ݛ��k_��ȭ/ 2��BdP�Â��`m�	#��� dyFeA8ap'77�����g��&��x�"�7ؠ����e�9ZN]�"�:�)g�A��+1��h�`oѻ�?(HǮ�邱
�^A8u��5"�Cx$��]��xv-<�=L�ʇE1��'Q�W��e'�AW!�|&H�l�C���W��˙��)9�L
A��lqAX���-s|��(��)����'$d	���E�S!���)�4�q���u�r��o&��BZ��XlxVHYEB    4f62     b50v�s@*1�����/�nt���L�������*޶��j�Q�l�.��XC�#�uN{��T�d���׍�\�q�q�������3ͨ�e�c��朥UߧT�j���X���3]�)�[Ս�<k1Q���ݗ�
�q4��[I={�[�x+�W#��WQ�G�7��]�{�L!�J}���T��	8��E�p�T�v��pȞ�`��#��4�� ��a\��/Utm����1���0�j�Ĩxe��?��{�����Y��^ F���7������7j��j�_ͪt�P\MY��T�"~����a���Yǻ�%��~�zV$9_�������2����1L�R�]"�*�5_���kʆX.����A�J����ls��>��@�D��f[=��R|.j%�0M\������ڪ)4�*�mذ���T���o�i�]b2�k�{*x1�ܡk�=w���:�iR|� 4m� ��M��rw�sD���$^MfS�X���s?+ku�q�aqF� !��(��/
y����x���O9���{2\�A��f��V��eƍ`욛��a��	��� �Hڬ��H�GǛ�Du��y'q�6x�3�S+˝�V�&��UXn�q���<�-��HK0�,��/O��吟�*(����ݪ��~^>iC�यܲK�#e�i$�"iL�|�vB��㼴��Tñ���#�|��_Z;�����ID�z�'zf�T�y�NNMVx��>�f�,�����r6>Yt1��&e��&z��>�s+:�����Z����P�r�*�4�K�N���@[��Qj��4�!r�N�B�c���:���.22s͎4��^��!��q���-#�G<�˗����}v^�i��cF�}*����sb
~Z{m(㇓.p���=�D�[`P����G�=� ���¦�Yk/|VjA 6��½u�q�J F��C-��=�����K�e#	DD�=uU9�TE��a�^4��A-ҹT� -�.�F
���A�&�9����O��V=Nmd��ֹy�A �UM-�"%*�i�����h��t�O"�oc���^Ẏ1�֣󯛰d����<;�B�T&��E�1�3E�%;�������3��kJb%����]S-��20�\��e�U04��Y	�\�ݑ;I��X�Ƴ%�+ɤ�����*�����[֐�%C#/펊R����'[ז��� ��S�E�C�wJn�L�ٶ&�$�E��B"ݙ�v����i�^�R�OѴ,O�`��Q�*�)o�42�{��s�o�y@��2�s��Ճ�U0���ؔR���U`9�� 8a���B��i��u" ��Ma���a��/rE������1mT%-�[��������XyT]TZg`*�͹N�6#����mr6E	�SM?g�X��k*Wl9�/+UF����%}��u܃����=#��A�j
9�^���F�b>����W�o	�AK/ӓ�ɪY�WO��и����%�+u3J(��:,ml��l�Ħ?��Y�TF��X["���I|�L/#"9hyZf��.�Ǉ��x��V+�T�
��>�=���1#�渆�/9��AV����:H�Ѥ��M�qG��� �֬l�<�7��ą��E\d�|a0٠��,szD5<z?�D��L5�ɍ�H^ԋWT��A%�w�M��s���>�.�m��C�P�zLPm�V&���4�O[VQ��aVǀ��"��{u2ꉓ�N��SR���=o���S<����eq�-� |JSκ��������8��%��e�]�=Z�}F;����zT����	�R�<��I�R�lw @
噴����ۉ��;�@4n�
ٲу΀^��x՞f�R��`e|� ������(��x4�MX����K��f�,��2��W�󈀬�w+�&\�=w��sb��& �պ�
����!�S�N�Z@�PFUx��.�tt�; B�WI	�E9����f͏���3��<�Nim�hg�Ps��2�,������R��#��<i�9NG��:��Gk��>�ӌ�f�2�ԥ��z[F�5<�����lrT�4; 2$<�_��
*=��!���t�q�bhК�B%��)l�AJQ�سyS��䘰�pUp��!Yg��p�T�&�I��*V��G���ɫ��xQi ���0�c�\b��@���"���[�Gv�fހ��ɪ���,j�GNF��\�G�&i�����q��`0v�{�,�y�>���;�^�x�����V�5'p?��l$��E�K�����L-`��r����
�@]�� ��I�L�Y�y�:�Lw�>��--�N���?4/��nZ�9�4�N}�������:��k�?��,�h	�C0{"Jb��#�dANVvD��3߬`���
{��V��X0�o^ǋ����p�` �=ݓ�����@�sW�W1����y�h�=���Ue��L� K<|^���2y�j�>�A1�Vd�A�����H=�H]`6VsP����(k\��$B#ۤ7�G�,�`[�����TS 7��x�H�(׌�=�R����l��?���dF�[5Y�5����Ҝ~��>L@x�P;�K�P	��2V{�T%�~�Ekէu�_��`�����[I�MW�$N���)4��cve�Cf�k��'a��v��&�ׂV;�E�plE5e&
:gN	���|gW�G��(t!��/O�l{�^Gu��"��u˯� �K"�Ǖ���&c/F�0qE[�	��U�W1+&bݲ�Q��D�w�`X����6�+XE}@�IϾ���l�+9�k���+�O�a�4�<�
x��#Ʌ�`��Ͻ7�8Nh�,D6���?H��T�e���@u� :���