XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Ed�:���++�?�.ˆ~��<G~���$Th�N�7�s���#v�"x��
�uQm^��GVSKU %�^5�,7W�?g�1��vØ�;U�#sV�q�����{��d���G�t��x¤������1�rK�9�(���"I��L�sހ�'����u���"g���g].?����G��6г�(�gt�`�B)s�M�j��fQ�Za�vք�a������K���5?�P!������i��^[�m�Y�0;ye9��6�f�|]��c��S2������\��r)[��Ɂ=���Q��:�W�y�K!���SZ%wgO5����~2�� �����/Z-���&��_���{�Z�8D�q+�N�	��O�u�d6T�*�#���|��i�'��;	WoC��o$C�JX�N	v��|�g�F�񉏭�^Y���"8�J ���������x�h����4X��6�},��DT֫���=l�2�l�mP�ht��e�G�`#W���3�CFڲ  ��@al���E�z�:��9,iE��J%E3Z�n�9�M�&u_���d����2�����Gc����?���xk�>ζ��e)��v�QQ2��5�m$7�cF[^46����yz��4� x��������@�π����)���j���FY�;��T�\��_1PG8�+H�i��XH�!0�1U��!?v�7��t��ț:����$)a����ܛ�JKu��F��52u�c�Ey���ml����@a�[V�)HB%vO�XlxVHYEB    b3c6    25b0�EԼ�!A=�!�m�mU,֞d0�_9����O�y��YbD%��A���Q��!4�&Σ"2��;�jq���6]��eUĬ�����֪W%���E��ѝ���?��r��׺>E}���0v�d�EY7b������W��o1=����O^-�S�����a�2_��Ԭ�;�5�X�q�BA���`mU>>��ܹ4�
4�c�Gp2{\�J/Uؠ-�
����Y=�s�p&�f��{�2�K��$��^ (��%�F��鄠�Ǵ[����A�l6"�[���Rz��*�w�V���6����^uq7�I�:���'��݀�h��3�jw�ހF��@~�bٯ�������n�#�C����[�����2�a=�3�<Fh�&~B�"{�U
$���޹��uؗ$��.��u�!v�{(kph�3F��&4�[��eR
���>�N]�K)BQ2 ?R�� 1�҆|U�`
I�j��y��Qfv�GkB7,����F;)&}l�$��C~	#ȴ]��ݟ�}�/����3�_�6������'�=�:��g5���$)����3�K	�u|��%�_l{����L���y�Q-c)�q7nA?VRC�^0#����+�r��LY�B0FI�fX07��ڰ�v5��^B�?�q~5����e�p�S��}7�JS7�S�^�ۙ����+���ۺ�nq=��$�8O�*B����_��r����&8��5�N� ����0�`ύ��aD��gb=�݊P1b�2M:�5t1Wx�wnVe�H;y] �GH���7���P|0��+�����v��Kl�ru�ֳ.������gp/�P[(�!"��ܙ��Ȃ���+�,Ŵ/�%��x��o���z���W%d�3�A:�I�&��}�w1���tz���ƖF�"5ʂ���l�m�����o^� 5�X���7
>+z��,T���=~���C�&/f��EmZ�"���x���o��x����+�VkD��A���׃�H�_tƠ(�"�LT}�kĿY������|	}k�Q��1YJ�߶�O	�����O:T�fM~oس���q>@��G�^ʲ��y��Tͽ(�����|f �*��͚Z��-�\7_���-��Z&�z!xW�,kw ����eL�u<��|��Wt,$��q�2P�}��]�oo�*�c���_`�2EБ�����m��WM��S�C|'�"�Ԟs3f]��:_�.���j�l)��J$���=#�~�]3��E��>�@o��c�|��7����W�N1н��6*&(����OL&��.�#R|�D7�C�O���(H����1�*�q4`���� �	zL����S�sQ���a���"2S��Dr�E��z�z$��W&�V����m�n��Q��ү4���j�ΚrpT�*���WK��?�/���8͌E�M�<��=�r}޾V�>�ɺ��c=�h��D���
.s�-�P`����}:���Z�< �!�Q/�ᣭ�_�X�)�ZR�����L���D.ؒ،C7�����.9�
Y���Q���'񇚪��Ƭr�kd�������5ml	�c�ɽSc����j�W��Y��I?��.	k���;�E��8�hg00nbH�'�NRS�3�&���P����V�����UC��kF����E��Ӆ�� ������� �v�@蚨�:r���Xz��c�}�{���S�P?����q��n�eԑ`��I�IK�[��s�k���i��F��TǺ�mJ��{ CbA���J��`PYd�웾���ڏ5���v��טݣ���9�.����1;�l&~�Z��>��f߈��N����O_ka]t;�n�oq�#��ˣ*�X?��[ ����P��L���'m����*j�;��÷>�u�7?_x\����u�����z���Y�����ӳ۫�s��u�;�v��\>ր����˽���P�sM�M�P���tǵ�3e����Y����_|��0��o�D� ���(e��E'S�L����<3�k1a��{�F��[�!��{��0\���f��@��H��!T���q�}�,�/{ؙu�X#��|�(h����rP�����~C����&��V�-1���Nt��������"�q���RF�fo��PI�i�-ᮯ�ִ&��M�[�1#�ސ�|Yg�^����ˢ#�Xc�U�On���	2��+J��oo�o/1���W�Q0���^!%�4�E���]�l��E�nB�JʹxĴ{ga�P�``��<ƞ��U�#���\�m�G_��	�6�������LENQ�)8�8�0����a��fp�9��!��,2}�Ƴ_��%C+�Ʒ�)2�[�g6�݋��i��S+�u�^����Z9���H�W�D���XⰰJq=V���������>}hw#�����.H��[�y��fe~}͙���=��w�k�u�t"�o+-[��sn�<<<-���?�wg�L����:�Mgw"��xVD��⁝Ɋ��r�DO_����B�]�`b���q�?�EuġҸ������[�7��:��ͳ��Ŏ:4+����m�Tt�
�V1b_�ݪ  G��w�$p����wk^�W�
��x�yAr�=pʏZ�%ꁕR�%0�P�Z1i�$��ҍ���o4%���o�Ժp��XmRjQEC��f��e�L�۫T>[�����!��T?G�lp�Mo���uV2)*d�� ��F�|T$�eM<M)�F��!�N.��r���d�%���'5��)ߤ�jn�� ���G"�}R�J����8��+�^P�_�^��~��*�u�z�3{T�d��A~q�XS�?!\B���x\�\D��rK��;U4.�_�`�e�A�*���p�X3���� ��������0������˧.0�ײ:�_v�X�\��f%�4,�Y\192@��ZV�v�8g���nTI^l1��ēc��3xM����NZ>�5��e)~9Y�Pe9&�],�"+��y0��s��Kv	�����ʍ��w�ԫ��l�:�[�s��A�e�_��U�Kt�_5tW�׶?\#�Á���B$��Ĳ{�y�U�I�L(]cDě<?�8$�����kp����
y��*�6���j�g�� !�>QGӦ$)&��K��ά�"ҥ��\�]/�b��P�3��na[��@A��iX���BG�R�\B	s��Be@%��?��)'B7��p6,�D�!�V��'*t��5���6��� ��B�=§�9vʁL�1�侓��I�:I�$\��_q���"�w��+j^ ��F�4ÌIb���P�L��1nq��络�>�!o����%!xmM��9C��Ը͛�ۺr$_y��/99羪�t� !R�]?���<�Y2�7�RC?k�,4����}��1�n��CH�C/��V�!'�ib�W.��K�W��-K�Z��~tu��0���aY��יK��N�����$3���ç��ѡ��zLG�1�yW��Jv2X`��K��b;.���^u��(�ۿc�Ӗ�p0�ݭ�^SIu�"D�P���
ul@�{p��>2����a�-o�h�dH���� L�hG�D�������qI���r�X����.��C9	����4����aMˑ�X��ʱ�y�E����]��@t��T�YK5���Р7�#x)q�)�]�)�.p�ssA�qH,aೈX��'���.юwNtR��-�ˤN��"�[J�E���;����>t���1���EF:���N��,t<��� Ԯ���-h	����=��mc(�ȳ�@�U�4S� �-��z��ng�C�╉S>LIu�Y����0�,�Z:����������mn␉n�2?Gf���6��5\������Z����I)<�Ȕ�9�x�]o)���q����ixd�U���q���.�Nh?j��xCDF�zow�a�;��:��O?�Pfd��%��j����7��Z�K�Y(7Y'޶cڵ�PƉƢJ��{��`c�u4��ζ%�U(# t�OLV�d��뼫
y�R�����9kl�!�a�fi¹Qq�/�ٛ��/3?�,@�=B_��h�1��w�T���¼��8���N�L':�c��zmIڃ�F:�G�� U/J[���߇����w1�n&�����C��2Oj��#��p����|}Rz�IC�Ҟ�I.��7��~T5,��4�f�]|��O|�L�~<+nl��K�����;أ��/�V��z��3���8�o:�!T�G��#=~�ޝft�� �w�ex�&#!������JZK�܂��O]Q�|���7� u�P���ϖ,�H���9v�{v#�tH��+�rJkfQ:��$n�Ջ��n�BnT��j���j��=J�) �F �37�`F�MR�-t�dG�0���]�J�����-�4���Dçf��P�W��3nkƌT�N��xТo�+F�;Ȑ)�R&!�)d����\���u}ޙi+r�X+`̪ի~�;���,�Q͊<~�=�eQ6Ô�Tr�ΐ�Q��A�G�^�wGF��gX�?�Ba(��	��&��p��T �<��h��	�9���;K��0����O^�$�;'.�ר�c����!��@������^�)4��f�j��_��%5�����!ׂ�atǔ[��MQ����uҕM�Sn����j yO}t���%l�#�ə�f4+	��_���{�/�0�E"�a���ńs��6�8�]c�5P��HT�@���!���_E���
���>� ZG�/�+mQЕ�9R��k�$��a5v�S�sfw�k~k�Fp�w�=�@d�'���nu=�qIB-�����X��c4�P
\����tT�Q��*[�)m�k�X7�YpR���L0�`�:�d������9JiK,;�Ҁǳd�M�A*Z�Ǧ��KR�΢��.;�Ϝ�M�!f[����'f��*��;��s\����*����%�<\{��+6��es��(zk17�xz=Y�����Zoh3��4BL�W�BkU��D\��cHY��%q����ג�����U��Z�9�ԛ�x�A+�G�
K���K�x��b�LI��|Y��x� �ьg:�\q��֞=�Q���L)a��%��ʝ������Qg�FpG��w������e�N��z��;��@�ӖZe�p�$��Ū&��eހ�}��޲�˝yb����ZyV�U
���u����M�3���Nz��d���Ɠ�u��Kt��W�#n���3e�GC�Aq����V @p����A�T�Z`�8�ڋk��Pt��Y��M]�WZί�'��ԠB�_�M]�GT��
f��� n���vV^\+����8@u_t����<Mu�ʂl%�-#h��x�[6=ih~6��CM�*�;�X4v���i��Bb�]����������~��1VMF�ԑ=��>19�5���,;�3-�U+?S�EG�n���p�f	���;�C���֖�|���c�jC# ���}2��q�Q����(n�9��>���!!�+3�����Zm����Ⱥ{� �l���SaI����Qׁ;��옷��݅�7S�Ua'����A�/�,�*6���g��E+"������$��a`�f�V�H�h�������*��S�� ����2��=�R���w�p�F���4��v:��Zir��p$MJ��ς�
�3�,�@y��={Sg�T�ʇ1zQD0������zLk_�r�Q�)���{N��p�G����J���Ƨo,q<�2�2#�t:3�"��+N&�Cڷ`�j-pu�B���f����
�b� �n�O�����~Յ��1K��+*��^�%���P-��.ߘ�H���$���&X����~�E��{8Y>=�?{��>Tͣ�	z�U��D���StP�����ˌ*���fb�K{{`�r��zh�k.�}(T���<�\Fi�a`S�X�y�Q.1P0K
�_�[�n�g� �����!7ҷ�ɓ�1Oe�KHg)�_�6�ZA�}���<U��6��A�wKnqҋ����3���%��Ì>�d�u�U4eٟ���o^oE����(�������qS�)'�g�R�����]�a\R�Wm����1&�"LfA���+΃��U}�d⥫�ofZ�n�"~���l�7n�Sh1`p��wQ�2�����/@M(��4:.s*����XL�=�I@Ğ�����dA��`�a�.�$R� ������`��)b9��=M,[����u��44mSS �le����<}K��@UI'fH�t(�xܑP��&+:s젪�s��%�OX:�)M��y�G
���y*q�ޫ�����\�$M��i$��@�*���ʝ�T��4)�n5��sv5�����6���czaɵ�T�X�2���WϿ��^�C�7~/�"�H����(q���`H�N����4M+���S��܃���e u��/h�>�C���@����S�w�'.�Z^8��D9ך�9�"�kz�]�~�)���\i�D�k[����٤�v8����*p�HY��t�S�h����2�,��d��G���E#!�W6w�����e#ڞ9�w�>}kl��s-����4E�~�&��e��F��o&�e��9�@�5��7�0}���w �ev�f�	�C�D����̼���˞u�h���#��᩷��G�n>O��7����ij����Z�<�;����ڧɪh2�U��b?��6�߸9�����	�d�d�ET�}�ю��'3լY��_�O�A2&�vc�4;6M�ͱ�;�f�������J%1���q.��w�?�&�M�v%`������r�������@v�/4�F�A&1�n��5Q�<E\,;���_�&"��Ozz%qF&y��`>]_ڜ�#�ڒ�ȓ5���Y����	����F�5�<�� 
ʻ�}��f�q�yD����Q/���_�Ȟ=W��)��W,���q���cU@�Z�	�s�ܢ/�$7*��u�}��ė4��T%L��R)3cN�#ח��%`m�KW���ُv�Œ��{g�D��ɏ��EeM��P;D �n�XMݤ�lR�AO�Y7�&�0 �0⾟N0���ż���aT���2������T*�fp�ػ�bG?�1���o��} ����F����o`��R� K�>�;�6�A�ؠ��X2!4���ؼ�E�	��F��F%�v�Ȑ;�����Rx���讋��(��M� ݿI��J�C��65r\��_`�@�9�ĈP���oe{!����G((�ԆF�D/���/��ح�s�J�|�+dᔦBN���J���ZeаC�ֺ�:?.���S�f����qz,���Q�:���>~��8�3������r*Qƌ��)�@�zt0oi�c��	�DU��pO�����N�e��;Eu͸�A���خL!���pW\_��V�˾�k�,%X���9�?��p�
!p��=.���A<�<X'J��0n*�AL`���2N���*�K�H�<}�ê&e�����	��s��m�t�xE4~�M����vJ2f��F��qup�;�y���}{B�>a��fd:<�S1)65���R�%9
�C�8�v�׳�~�k������H�5tYYPm&� ��;Z�K~��U�ғ:��AݓBw�ukU���qEx 7w�6�L����K(�i\��I?j��v�XR@X�O�����tg6i`�
�Mr���'U)Ķ-��G�m�5�ᤥ�Ē6�2�XB:�����W��*7]x��XQ�����i��[��Iβ5%�f�Ay�ϣ3e�VrM�*�E;;�q�Y��U�Y���m}���dx�k�xc��@J �Xz��|�DSG.��b��
��ˡ�\"��?���~��i����� h�	i��8;=�Q��JO%�����+��)%Q�h1uZ�F��Lύ$!WU�E��G�?T�a|l9����l�t�ܑֵ���:�j�AD��F��g�W����+�&�����6�g��'�n�}�Q��B���w ��?�1������ �lx��d�,� m ��R�`�&�� �����oG5�GvU���<r��Z��
�ܠ昛�e`�O�c����Sb'�q��s�����Q��s�t%��Y�@��QX�CD8������7�ѱU-	��V"���<� V�ũU;пQX�QMB����G�ũ��-|�u��l���_�����z�k���C�l߲9���!�{}��Q~҄ �Ku�.�]ew���T����A��dOl�[�9FS�4�F�]�B�i$Ny;Nv��L����Q����.V���<� �8UR�V����>Ǳ���?ykT���QD	k;��Q L�K�� �������iD��89 �vnm��t���0�7d��2V������Yv�>gOd���vL�D{�,����6V�U���w�����p�,�F�cP�̢>�ޜߣ������A�;��{u�s�|�J��R��@�l:��� u;��OXX�>��ld �p�>�1��z���L���p;�C��1�x�S�������9��|C�N������3�m�X +��a�5$���h������n�zI�����T��{����I�M��Ƙ�$/�EM ������U��I����a�5탄U��|Ҩ�������>��5(�Ĳ�z?�s�L;Y����=@nU��	a�~����r#7\,,N����4uCR���T����<���ՅHq�CC�-���~c�l�XJV��T�p��BK$q�X�
�,�L%ԢP�X��Zˍ��Em&W���oh�y�8DQ؅@��k�@�U��}�S{D�q�g�%*[�Q~J���-☲B�oHf�R$9���ɼJ�5�~3�4���N��#��>`&
��	%��@�tݕ>3�/kͶE�t�\3-�A��~�L��:�	nJ�M'�dN훅7�Y�m_��׆��-}6�{:����D�_�5肋1�����k-ȿ2��6�x'�Q��Ď��c�e�s��;^ddE�b�S��2���F=`��ܵ�P<£�'�e���
4������)��������}�d�%X���PA�1._*�$�\<��a��S���@ygᚹ!�Dޘ!<pg��tU����K�(�j5�K��c��f���|B��ٍ�w�+��8�ŕ�&ר���u�݊(H�M�\8�Q�
�MX[o�k��s�Vɬo�f���� �S{���m>�����i���р��I$��_�,fh�L�	5A�:�yϷG�yO����A��[��MQ(�<�� ��k�W��؃D��*�lZ���޹�6���2��1��Zk)C��H���'f4���P�2����7&�C��<-#�9c�	��->R�-�LQA:�BI�C�P�ԓ@��x��>�' 6��w;�b´�t��s�?0Q�M��i�b�&�j�!Y�2s6���;��^*�IzǼ�n+R���pF|��+w	:>2�0-�-��eK��