XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����="Nt�p���xG�m�ܡA~Qu6�jI/|·=�bޭ3�`��ʃ���JZI)�q[���>T����^O��{w�%���U�Jg�o�h��i�Y���3�ʕ�Fa�j��k�d&�F�(<}|8��_c���N�^:�Qbx��8B�d	Q��x{6�Ҽ�]�L��o��ny���6��eK�񸏘��Y\LH��.�Y�K"�]F���w�U��qv�-�d�q5��3�����s|�T���wq�_�se�c�x�MV].쮐����O�L��ʱ va3��6"c#=v�!�I�@�%��/����6��ϰ�ϢK$FUŬqu�HO25�k%rO�F;Na���a�����t��dsk<�a� �X���C����Qlw��6f�i�8��\�Vӝt��s���P_m�#��8�;�/s�`��F��/�0�x�YKHnҠ�$!&�� Sv��nu$�-ן��aK�a�`�K�8ߙ���/.v
����sۭ��7U��ٙf�Q�GJ�v>�%�o�s�o�/�3�9�DͿ�m�8N��ԍ��4�)�@V�T����y(k��VJ7�
����*yQ�`�Wh-��;S���zV����ނ�W�������Wy��?��r���JB�9&D���]%�Q�`�񣀩���]��tzi�l�1���f��[a�Ns�������1怱$�>u�V颦��.i�h6f����62tgk.�dür��#��7�����Ht��cN=�=t�'�zDG��X�s�XlxVHYEB    6346    1790d�>Ӱ�縴(�Nu�X;v6{Q�+� �荄�`��v0�����մ-5gǯ�c����]�����f��5�Ѭ4-ꗑ�2�^���B�ܙ���*�#?)�yé�$�<5�rz��Cﭧp@�EL�M2��}6F7��dņpI|�T;�5N��a`w�"V΄����:q�y��N3_�8�m���M�(@�'����W�_m ��D�ޱ�L�0ױe��T*خ:����[��D��tbR��N+k�� l���x��.2׻A�%��oz�î(u�a���ȶM��a� ��8�K��V7�v�%�Bd��Q�֍;����{"�h�>V@��K|�
������h2Ag(�~�!P�Ð�����t|vi`�V(y.��[6,��MM���y�LR0�V ����*7����oQ\�����5���$ڔ(x�����7?]1�ǟ��[s�Q�A4~v.��}�U�L/n�72#�����x���}��O�Tr��:�H�ͼ| �l�� o'�Ѥ`0�i�t�X7�uB������@�(.���������|�)��������>��"%C�GW��.fu�B��s4�3��/���l31�MY��
�����:�^��g��qVf������և��<��e8��1�Q)�#Jd�, ^������W՝�~t[iJv�#1_pf=�o����1-���CbU�#��>(*&�oh�b!��pv���ҿ֡�dEix/�6�@V5M`Tl4o�[x��K�RS[#B�}kg�q�a�K�b4�D7C�7U�����	���.u�`�y3oR��|�V8a燃+�8���[�K����R;B�Sf�R9I��Au�͕z[��4����:C��:���5<�6����|�4�8U���N��7ǳ��񍻫xM�`�5).�����k]D��w���W��'��3�o�qv�5�v���ڪt;f8yu�`��y��SER�Ë {�u��(G�b��O�6���p�P����[��6cˎ�U��էn��q�2"��5�;���9"�@>�%M�y3$ׇiz^b��JXw�;u��TN| @e��/[@P� ����>��j�I7AU��ZO�\�Ŀ
�Քi:d^0�]��(��R`D'�-c�NhE@L�04i0öE	�̟���)u��g״�,.����a5
ݽc��^X#g�`��wT���j/�2�8�dM6��r��	G�/��(K����g�x�w#؝;Ң�[,��z߬}��4�g�꒞���m%2�~�E��{~�tv�-����.�om�5J���۝�4��l䵺�g"<�6��:����������������l�q�s��O�z6���mPV���y�ev���c���߭��8M���BZ��n!�s]�Q]�	�=ڔ�\t8�ɦ.!?��cm���g��[f���a8�;�N��͋¡{� �
�y���Jl�6o0�QB�� 7mi�a~�3fAE!�=�J�?��|�l�9jA?n��8>���ϣ|`���F�cI��ۢ".A����*M5�'�	�L�!24t��I���j�"w���;���_DOt��W<�� TJv(-
�a�f!���?FH��Q.��
�2���"�.�z��@���a��"����%ڲ�KQ8'�v�9^z��~�
z1��?1�,�vi]���vP���X���mIG��1n��@kS�W6;�iR���F҆��a�0�x\�\���ϧ��	9�H=Z�69��د��H���e��d(��\e�ܵ%H1�Kc�sC��v����XT���|�Oha���,���rm�q�%I�fW��MA��I�L��P�����+)��UX�`eHo��P�?�B���?m����-uv��*��b��CE��w�*�Љ�-.��M�|�f`YjP��a+���Uyhh��Ԍ��ųx�jy���J�Tհt~������%aA�գ��E�d{��9R��e|�|�٪/®M����p����|�З���\�,���D�	��������1:����s�'�݇?p�9$<���^�,��ceU�KX(�AAã9�������ίY�W�5�%�'�L2WB��`����]��i�}�H�˚T������3��\9�5�y~�'ػ��::_O�s�V\�~����$j>�7�+/�E��#;���Z�j�+M_+��3ص�B��ɥ"�N�.w�jIb�*[ �QPR$S��CYJ�XN9���)���Ё������Ԩ���!�g��bue�g��-c���9-�/������|�R���ۗ�ƫ��?������-��	�|����ǒ��V��.Eb����O{�6Ɂ��g��b��¹�l�&�op�$��l2B����m�M���.�{PCn��ب
&��ĵ�X11���c�'���PK���
�����0��E�b�<"��"}!�������x��4���*]#xj��q���@^&��9)Y_��I�,����*���&Щ���,��#�;�PcW�R���Kgi�� �>��N���>�ŧs8��;��
�Z��3�/"�4����������}W��ĺ1Q�E⧕��v��r�V������ ܽ�:N�1���;ɣ0ʻr6N|�@2�,O7�	K�%ga���XrU*�~&��5�.}��NJ�F�����9�Z�^�(�{Y�+�mb��L�U�=�7%���x�+�C�\��HVY�Y�\�X·��-���QM�:ž�0�����_�������P��>K���!��6
4�m��njq���Pt�_�z��$�uW�9wH�����_	/r�Z�e1S߶zJ.3�"�cl�fN)[���ᴚ���;�u��AWW9�9S�!��>£#A�������&�;I_+L�6o&�r�$�T"Z��ƹQ�.������"�M�I�̣�h�qD��R������j��3�'1�v�`�>ڄx�s9oǳ��³��T��h��!�/���M׻�X��.z4���i�[pn"'Rw�PPI^,�!�,� �?	f��M���2a�Kw�Ѳ�����`��8�^������G�9�j�ڂ�]�[�3q��q�;��-��Gэ�uɮժ��fE��@��-gno�w+¶��}}�K~ij�I�f������v�ݺ"�U��t��� A��e���FJD��L�)-ƃ�-
�(��m0�j�	)���)}��XTRTk�(*Q�i�+�䃩��y���7��+Km��?7�@�\�ZYJ���A��A��g��NG+q���#"�m�S�g����_S�a�����V@��A�l���_�T5�䐋Q&�j�Bi�!N	��u`��i�{pO+02����>Ut��#^� �Pڇ"3LX�!��>�z(�Ј�w�r4����Pe�Z'Ȃ����$Sf!����ŹXx�=:m�����f�"*+��H�lM�xh�p�+B�g�KV*а_���A=\<���)ӴA��vw;E.Y���lƚx������<�K_�^Q�k��.ޛ��f
G!7 �%�\�V���1�����J+�*2`+1^���M������U:��J��#����sC�]%�������{燻��U�2�6��@�Ѵ��O:p��zܑ��[�;H5+g�d���5�p	�}�,Z���[�����.��h��K��=Z]e���k�?4-^�"�5��+F-/�-o���߈1U�cd�y5��d�">����*�yR����;�q�d1t�#���a��~s�H���񪃢-C+�������C��9x�����iKb/ ��RM�88�q)`y���>� ��I^o*��V�3�LI��Z���#�ȑ;*�|;�o!������6~�bd�p���Q�󈃢	+����0�Ut��IYwz�O��+�	s��ڎC���,C�˕����JAP���H�������)�|���&��)���5>f�f���v��͑u$�12'n·/����r���f��$0����Y5�r�p%/%���e��m�Eܒ[E�X^7�?��P"椆��bz�������ӡ��u�����c߼�j80 ��}�N��������ڐZ�JnP�yV��n��X��lu�d�1Q<��
蘤�)���'t.&;�zC�������G�͌T��c���̟_E�q�3;�x���Z��R,��כ �BuU_�B�x�e A�� ��� =E���\=X�>w*�4��X�~��E� �����Մ��1DK��:«)sR8I���TZ<��C�3�]2��lMr��G(������ ��F3$�e}�Y��;�/�"������>[�/F�U��XЀ6�lG��Vj���f�cF)�b�2�Ҵ��}A!u�/��:c�e�y�����U�>��{(RS}��?x[q&e���s�j(A�z�;t%H���;P���"�JQ<gJ���
��2`���/���l��X��y����c�`}*w�z�iG6���|C���Э�~�6�>�$�+�a|�q`|������Z�Lol�CW�1��6m�S��6�<[A�򩕼�S���%g<��i��[\���\S��� |��4��}FF���*ߋwC�e��� �-��n���f$���
 7��&�fw��C�� Գ�������ҵ)k�d����gϢ�nh.����-�zv5�#�^�3�V/r|�ڇ޳�
��aW,9#}�ؐ����O>��L|ڊ�\��Q�N4���{���Wi|�Ai �f�&��� Zw�2/m��Y9@ �E5�qc�R��[��F^�✎+�tva�	�X|ɨ�yr�g�}�}�K~�F&�H�F���F���H�BBf�q���K"���8/�Nz�*fڄ� 6dt�j������$��"�����TGoړ��Ys2��8��r�5��8��@�ғ�4G��q�����1h�g%��t�NO��`I�
������s��M�4��~H[SN`pB9M�}�Tj���>��["|'$dR�)ڳ�� �7�`E�QO��;�ԏa95�����sg����X[=����H���qr[� *��C�4
�'�`�8.3"H��qUN������G/F�[��"�s���2�f�(C�WȞ�ɘaT��@��P���D�M��Γ=	��z��q�0��.
���ӌ��X#n���.�?j�Gho��V�'��HFWg�-�X�����L�H�PR"��8�)�����0�=,��T(��c����b��y3��,[���C���^+���Ϗ�t��H�˜���Ð����M����N1�h�͇���b	�w���9wĮ�A�i������o�䙬�p0�!4)��֕M��O$�&�b?��6�C�o2J��=}�y�+�gKҠ�_^|���֓�� ��#��+�J$Xu�-���r�X6���|m��y\i��� L|�u�������Y��yv��vw��w%�^��`m��iV��=���2���D��;��s������u�lS�.�~%c�xZy��L0Vj$�b�MR��,���)��I9_1��ٮD1&o���꫖?��4Y5�|9в����Y�ƓZ��?O�RaB�ۉ���c]zʓ{�{&sa�畝dk��$;d�����a�d'��M�8-��y�P,�ʷ��'-n�� C��6�?���G�#�u����`�,�q?�l�"O�4�m�җZ%/a�GK<w|+#��hHʫ��S>ޠ�!�����~���%'�Ő��i�䏏��侬Fٽ�w
���@~�Se��݁��d���?�-3�;�����̵I���1�m� �r����.��6MV��:����k�a�d� ؔ+�G�טL�*���`aOpj����\��Ҹ�QG��Xs�����xГ��h���'���8T�H����bW��ڽ���W3��8�#&�s=�E�&�['xS�V���?w����Q�I�ʷܱ