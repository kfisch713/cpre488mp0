XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?�� �n��y8yՅ"�C]�-�.=����˩x�j�g���9y��~z�m�W��ֆ�B�q���`#�܂c;�`_4�`��"t�hb������(��2��Ky��#~v1E�g7=����Ck�;�,�@M�Ɣv�si�a֪��f\�3:��g��AzϓEi-.����;J>n�mK��J��H�������n/���j�̔z�T���5̧.5ȫ����F�*�����g�擏tx�r-�]����e,�
���e�0�ݖ��$fgI��($�r
f�3jz��|��l� �a����l¢٨��fb��и���m]޹[W�a ���;�����R���Sߥ�#����R̭��Nsx%��"���d�T�t�s�� ����� ���lT��r��wN/@�CL�X��y�4�Z�()n��"��P�v�+�\{�*���n�ȃ��(�n��d_�ݻO"Z��]�v#eʁ@IU�z�fO��0&P�(����4�w邟c��C|���)��R�SM���F�'��U��o3o�H��?].�RҨ�\��I�e;�v�u	���E�m�,#y;��vPA�dG�~���q�RB�]�#��]�Z�L��UJ��<9_{:\W[��'�J�_A��vq�0��E{����3!�M��"/{��''G4( Q���X���R6��!��r#4i�nfzU��Q�T���w��L��ڔ�''���}5�����`�l���v%4Ъ0�
�C��z#^g�PXlxVHYEB    3fdc    1160����7@���w!Ȋ!q��9 �A�K���9���ʞL�{3� ����B3Y���{����w�\��^Z^iA�<:�������9M� ����$�]��K����h�����7I��E�e�<SsЊт�ݴ�A���컾�����UU��:���B�4��� ��G��ۇ08A�pT�O�'�57iQ}���1��R����@���h؜���=A�%���]j�gt��{����l[A���L�'�t������Q�qV���M��_]���M��T?*�:�i�_�i0��P��	���Z\o������/�ɢ�7���I;�8�ե�K��:nL ����s'ם@�{�K�S�`�1�n��h�p��:��ݸ�]�F�$ �Gm����4/��l��3pQ^O��K�oEb�Kd�����4�K��}o��I���mP� ��=���\�T�.�q�T��F��q�B������� �}�Z0n��Zr����0��.@X���%	��1%��ǡۊ����o�v��N��5S�gH�(�?����-�W��^�-�������b��B~t�5�ȋt,�Z݊[nϳ���*�=�T��P��?�T�?�
�8D��+>Յ�#I��s�띙q����@��7���[G�G���d��k�j�?0��� ���:�0u>:v�"H�U2莰��K"�x�؎
��s|ޚ����ذ�X�0�n��Ew�x$y$��YM���d�%z�>��`�ve�gĶz�� r<��y�� Xo���jbZ��?1�`dIj�J��:ݎ��JyAu�gw$�����}��-���G�d��Ь�v�2{|�d��?�n��5�/�������LA������7އ+���Kɨ>��z�֕��g��`��pں%5AY�7�3�?�8U-����Fgep�k�͒��`���O��>�'9���!�U�y.xq�#/���ϰ.�V@�"�������5����;�@<w�1��;Yi�����{N@pѹ��(��k�����93yӣ��#	#�����% ���7u��aR�����ء�ev�4�+���gG-[�^��B{h*K,�S��!ǑԮ*��\ T���U�n�聧�0���LA6�"ׇ�4-�Y�`��e?��x3U�����<�Өx��pTB�DB/���MA^)2����3>���,���s*ޜvx:���%Z�k�u�n�c�	x>�=�[4���y��~�����C�B����ߢ�m9�#y�=*�s28�d7�:��YX��H�~C����7�8M��1];�BXcI.JL*K��+�^K9���X���c��w�XKT35��}z��1�����۰p���x� ��~�hު}��ЊQ���y��*m¯*���9�O.f~$�6FGx�,Vڄ������o��g��PM�n�w5���\�5˥�'^e�2(�>6?ݜ���w޸v�񇀓��3��~/�R�_�̦V�C��d�)�A;�H���i)��1�%�Kd��!�u��o'�A�$FȞ_�� x�~R�` s<�(��"�\3�U���$z@h6�lo�x���~�ͣ��|<<G\V�����n�F2�ޙA��Î;�½ bM��~a����=��1(�b���3-���A�w���m43A�ή(U�)`�c��b�ntd�y�Rm{@#�Y����T�/��+/a	�GH�ZG-Fm�O��)�,�n�y\,��1�
��c��%��*��C��`?�}�W�F�J�w��fPh�?���]$K�n9�ݒ��2ձ+�<?��:�'���٪H�:��B��q�Aˏ�r�'��f*f�o,*{uS�jaes���F1�@ԎȺ�rj���s�l?�q��jQ�,�h����(5��c�7il5��N����{H�F >G��v�*�_k.�_�NFJ�N���-+�L���u��r.Cn!SG��M�C8�u|x-v ��ZBL����L??����F0��k�?��楢�'��S�2���5R�������ߒ?��|5892��h[�=�-�(��2�aʡ@w�X`��1�ȃ�%�7�fbW���A=�z�c
k页b�:�T�'�zb�j�IW-(M˖
r�.�I&�m�X����c��U��]��9���_m@�$���e�`�8�	3�8?:�{E����)$s� �r*^Cs�M/���=\����'c�R�YƶD��1�H��tm����o�������#˥��Ę��>�k-���4�J�4_%(���;f�l@m�~��#���5�����4�y�uw���R�ds�*l;���F�x�����Xm*�뾑;".�����l���2���d�0>�r���k��&�R*����1�x�����I�F�L�['�v���Tu�`>|l�}܃1a�#��c��k���l&H�;im|�z-��/�Y.,�,Z��ImA�wM��9﷾Ҙ����ҜIH"����EKΗ2��r%~��cioJ���/�i��;������zN�(<�M�Ł�C_�f�N��a"�?[�*�>z#I�7O3M@p�=E�Cݡ�^Ws_ࠃ�3�r��A����]�G�i�IB�4�"GXn�/w�6S�,��e�V����a�MQ"B�Cv4u=T{5.�SZ)I8bO�k}�L����~�ym�=�r@��nu��9�	j��}�#O϶w)�����<����p�c
�b8I�QN�3�E�
EE��a�m�n�-��ˢ@lV"M����|�(��Uf���Y>�����.�!�9�}챐6y��;3bx���ģ���UPn��*�*�L,`�)NB�J4�VRUßl�C�QbvЇ��E���pȃ���*R���q�W�A"}���~9���r���cA0��V�����8�w���k0_�����JEMy˩0j� �8�x�:��`myV�1d66��Ga�������"{kկ�a)zǗ����p���c
�m�ݕX�]����H�1��`�]��Wu\ݏ~�Q��&��U�7;!�U�F���:���Ʃ��
�����`�~�a�Ɍ�p�oS�` 0�������ky��!m<~#�A���..I��W��<�����!�Iqq_ ��@ٳ���;[,�#s�<�1�|�;��l6�8
�����	��J\���5$ ���
q��U�
���~��r�S��tH�DE1;�=5���P�&�'Y�Q�@m�w]y��/�;J�=���P(Bb�9E�j[)��c�$�e����1g쩽�h�ʜ��S=M*�GԂ��w��f-��c�55�}^�=�������/���u�J��4�Ξ�݁<��=U�|�y�.5���aM�f�ܝ�N=fˈJԨ��9h!��b�	�O���m{���6ɩ�>m��kL���i�~1h{9?���N7-Q�ẘ!�*9�G�Z�v?9�q�lp���w�5����ƻ�Gn#�.��R�*�*&��ߣ��]�XV���t�IkUS�J��2��Ju�8���#`��8���<"y����ٗ���N,���'oO���"$}0Y=.�v�e��
wF(�M^�|6g�D�f����A��Z�.���]jExA3�(6M�ڵaI!Z0��+��d�U��� ���!�d�"Y�e=���]-Z�9p%�f%h�F��������5殘���D��8�Xo[x�U�c�!!��mqYɯ��� ��:�>&SD\�=���t]�	�����~'@U(ɏx��=$��9/���(�n�kgt������c���'���0�AV&�|���AoG��fۂf,�X��^�C+�vgh�����:���e�)K����0�wJ;j����}y�&"��D$B<��R��A�|3�� x9���dݫ-u��?�mW���@'�f8_!��>˔kޡ�h��X��kg��սV���fboX�`d�:B�Y3�	r�ݳ�uBU0[O%�E}C��\@�-�/EtZ�����D���+,�����Ma�AhoMbv�%@��>�:�0�z�CM�"��j�F+��G� FY����Е��"̱�p��Ad>�L���I�$J�z��B.F&����?в�c��:ZAXhC桅ڂ<���R������xO�w�;�b�Sf�*� �u\3i1b*`�k��D�ۥ�p!�i7M�p:���c�^�g:��̓��|?��ޅ
c_�u�0j֢
�qw��<���z�� ST�ߠ�y�lT����#x�a�6�ᵱ�D���"l�W�'hj��'��N\KU���eȌ룠3w����������~�C�鄣��ˡ.{��2�4Z�}
j|	���
OWS�L��BS#w��7�J c'~ J��!k�lɔ����I�)��c̅h��vP�V/lh�\���P�puHw�~��؊޳v�⡃����y�?N��iZ