XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Է��Dv�t��	�V�ܨ�?�0]�	�2�s�޺�����3w==�pZE�|DS	z��zqm�Ѓ���]�d�л{\�>��J��9��Pz�^������]�N����GA�$G)���RLd�C׺��u��-#��l��,��a�	��&Ϝc�Oy���J�h��5t�t���[z!��Q��{f{�7�=֖}J\[�ඃͣ����t����l�|�41LR��^nq�`����#D*@;)߭m�e��-���d)l�.K0�D6O@����}��	���Y����aF�&��O�H�xy��`�g6�4lA�j�~ฒ��������^k�%��3���v����_V,�8�+x>3W�U��:ĄO-+c@Vb ����X[��ߪ*��[
���p�3t�"�xd$>�6X���˨�l�q�K8{:vPI�+/�g�,P�lه��L|=FW�,3����<5?4��'�jM�]-p�2�F��Jh���
Gme��I�%��E��E �����K�Ð��*�*.�t&m���$�,`�Ґ����l��WW�G�WuGu v�d������u��~���״�ˡ�h7Z����b�?*�
�KB�6��t�6K�.���@�Ϋ�@�͏?}Gx14&HT���n����;7�K����\pH˗'�|KY�^,[>t���)x�{sz�s���y����p���q+�D��>��!���X]���
�޿U)�<G˔��e��I��Pr*fx�	ɽ�K%��XlxVHYEB    b3c6    25b0����&"{��R4+���c#�uk����X�V��3�?b�x C��e�~���`������/g1{Xl/�cĚ/F�DT&�E3V�a�Hn���XT�������>N2о���ɜ�⫩�/�_�E0��3��0��h�;�#-��^�`qo�N��nY]�2깊}:�am��=�1f^�h�.������ f:HTVMKn��crp��M$KW��T���=y�]���� �}�h���!�#	��3� �f�$�����M9B`�ehf��4��7Ս&%"��y��Ep�W��3��L@!pr�v�����}N�(b>9QlU�r.������R�]0�i+F����[Qa6g��y-�,8���qw�m��y��u��fR�5�:7�~O���Xp\���΃m0���b�h�o���O]�GϜ��(���@`���pOk
�$?LQ�:Os��1���(����dH�M9���_��/	�ף@�<Y2
�|	�[A%��P�-��"#�b��R4��F����/n���^~��^l���-M�!���g�9��ͷ;2�ix=^1�K5]2�-�ϢNZ�`1���=衢6�3��c�!q��@�Ǐ�T\�!s�'�J�ڣ����v�B&,��B����	��4���y���B�����,HG�ϊl�d$�zr�L�z����B%�����)��GK�U�+�S�T
_�(�O��Ś�
�ѩ �����:en�\����C n$�����J!�J���"7���B:�����*Mm�ep�0
���VkY
$��V����Ғ ]Z��5-��-w���C>σ���Q߮X���_�Q�*�"F��$ޅ����A�Z(^�S�����UzT���m�еa,rc��B�֛�D�M�����[��^\1-;-���oƨ��ƞ�V&�	�{��T��XWi؊�Vi<�f�0E�8�4����XVAt��$+�꽅�$�X�!>�B���uK�/`P_���T��"g��p�$�� �<I��*�|v�m߰B�Wܞږ�$U�F��ac���������t�C��͂3v��c%�](e�@�E�8�!9c��ZH&is]dj?7�E�7�+ڬN��J��[�j.��d~�G&'_uJO�6�7�{�n��G<�SM�7B�N��u��Yd��I���0���[�`OI�r͒,BqXg�iR7�.�9�"y�*�vy��W�0GA�j�~H�mv?W�|�o��$r����T���s��V��э���_�4�	�yu�(�0��Ø<�¸���l]G�I��F^$�G�S��J7���\)�����'��_���}�b�o׵%���)�H㵐��W��` �����7i���I�.V�Fl��5Q�Q�Ig�j->�]8��*�?�B�).��n�[*^�gY���}"~��*,�5sB	���}C{k�!R�G��Ǻ0��Ӝ��Δ!Zj'4��`���j�[w�����{3H@�7����%a�z��R�j'�N�B��䚬4��?Y�1}��M*����Qg�����D���n��s`�m{��~0���Tc�_� p����hq:f�9�bG��M�kmv���rOΖ?'Fz�0RK��$�i�,À�`+�0æ>� �șh�"-��/q�� �?f�y�y�C�
vw%���-����.����)�ϊ��Ai���¨?��<F�e�sKR|�OZ 3�����������{,�z-!J�� 㳀I��U�N��,���Z��=r��:)�<b�CXf���v~��m����LY,����R������fy�r�m�����J�D�d:��}��8�+#�`/Ns��ٕ�(��6Z�D{aم�<�,��c/�z�}�z٥�N�1V��K�U��q�u�U�_ଠrC��m�p������n�=���B�8g|V�R�i��X��w ����r���*�)Ղ��Ůp \�k�>�8oC��ʥKqЁ<;�Q(-��y2�~Ch���7O��=��n��
v����H��$.�|V�OeQtdI�	7���I���N8��Y��"��t��Õ Q������:�����Qq��������1{�h���*��Q�Y�A�\�j�X��rj�o-q%�����B��N~sn��O���t��:3">�0������^ꕪ�Ə���"r�f<9ZD]\�w����vF������-��"d��=cP�����J=�L��堚��P��B�b��ɂ��of�����L+�	d �� #e��d���ׯ�Ʈ�P��dzԁdM-ϸڬ��G�D��:G�ŃDl�G.MW�~�O�� T�sGE�Z����y8e�;���v��ۜ���j��-8k�"�������R�W\��®���P�
bJ��2&7�ZRO��`s]��"�����)���׭ݨ&ua�+�-��|$�)n"'5$s��Y �}��N��TsÃĐ���4爋�s[&?`�i���# �P�5&y� ��o�:R��h>{�L�}"���R���:O���� ��L�P�;�Y�k��B(M	u^T<�Ii��dcg�&@4���y!���NH�\t�E��v,�t�`�_^����z�Ikփ��{��> 
�Ȳ�$8�7�����x�v�h	 ���0��@u�#��{�N½Ո�z�S{%h�8U�.��xr��$j���̔R��������n�q\X��{Cx^��)F�/>���8q�I}��H䡨�p���o	4p�����zGëhE�!��|l��Y^Q>ŏ P���G��۠S�$X"�7�e�O����us���@�ǆ��8c��s�g�Z�o(H|!
��:��u.R���Y ����]GUu�Cy���Ui�}����C�S�!���oUQ>�%[��P�Te:���)��d��e�俔e��
�]�z��gT^���{�	y�5uLN����1��4��>l� B���姆�G�Y�Q\��P�N�g�'��;�s�������ZS?�a+g�8�Y?�ʂ�̅��q�'z�୓c%x��L���Ev�8� ���)��Q>�N=�Q�a�&�B��&%۳-�*��7��c�
�|���p�@�h|+�M�@Ж^B�(A0�qx]��{�w��߇�ԑ\��s�3-���_z76I���j�������֌����/-�KQM-X{��.�,q�@:�(�;X�N���cdT!�46�t�йq��$�G��l���{�y8r���9���3~��yP��W�̯c:؄��8%��
�>ÝfM���9�?Y����)bFj%;�OS���A=A4��4[5��>���K/,�{!���rO��-�D&�v��Ȼ��N�4{ ��Z�gau�Tɵri���e����M�A&b���X���{+)�{�笅���[恻]�W�P�� F�8�H�eϺJB���]*]���JƂ�t?źU���Q�������q'��mrƎ��=�����&-��t4 f�"���B��ق]����s��f:�g�ą�����$3M��j����\J`�T���v�#�������2��ye��zܨ�^�ad����(I�0��d3#�ο�գ.R�����i��f��Q����&���/�<Z��
b����۔'�o�8��c)���ʫ{�oS}Z�ϧ�[��\�!w�X�d�u.zq�w���7v��dR��%Ѝ�Z%�#@�G1�]���	��c�A��<&��+vf��Ҍ,\ٗ��č��NV�Q�!�[{h�۱�R�_�� ��n������.�^��0�^iy�}��&8}���SVluSE���Y�Y��������u%�����/��L������p?�J��lN��`]�pL.��'�F��Z������щʊM�R*�g�Ƹͫ�]�Ϛ�S&�
ޣ��.�T�Gи�d���_�:ѩ�[�n�N\_������ۄ�d��5�hSNy��wJ_�i�רÅ!|���^��EA��+���F)�Ľbq��T<P?Ѧ��faC�W�pB�Px.�w��MUWrf�q�#%�C���m֊��k�:���|r
�T&�\(��!?�]��W4��-W��^�]q%�m����'�Q��0�C�paԧ �h9���ݞ��g�|َl@d��.g��.����tna$D/��,(�%h�Q���.%��1J�m�V���5#e� � N�d���bt�995�}�|@2��&�ڱ��Pn�x��;�f���� t��u��4G��`��_�v@:t1��$��zO�k�5ċ�0����٨�j.k��7Z9"����;�L���.�u%Mk!L�b�]��6�5b��m�$�����z��B�������Y?
����6S����]nP��{��zp�
C�H��sh_�eQ�
,�
s��	+W	��+�?�fG���(ڔ#v�H�EaS����T��Z�sd>�Qk�<"��YwI���j�/Y@�U�%Ҹ�v#�v��!쁇)���4�Z+���Ѧ7�/��~#�rb.�Q�/F��"�Q��_cݱ�p@��*�@����ԛy;��&t��*��(��%�����8~; ���$�[�W��W⠨����E
�1��>��	�-a����$�\Σ�I��SP1'�����֯��\�x�q\^�9��,�Y���Gt�����`��g��f�%@h��bw�}�v� TsJ�n��잿f�W��ur-��KO&s G��mg��){�Jw=|_qv��N1}r����V��啖���G�M_�R�ul��:h�6����)j�[f�r�2��^;��������J*|��s`��B�U���8y��C�k�s/l�o.I�S�n�l�)u&\ 6{{nKRa��9M�I��^�7��#,W��~����h�P49���g���?�5|'$��5���юJ#�>�Y�|�i��2�L|�C���]���u�D���}Z����D`'51�8��+��d��7�:��0X
<���/��=�����s�\=���f\��j_�#��{�+�oO֔��+��d>�XrT�7���>�.���ɻ�:��ܲ������y-z�J#8.M5�.�[Px��"��.?r���#`���$�˚��ˋyW�B7Z��%装.z���{��Ͳ]�9�[/u�O��bI����&C����<�p�FX;���0�r8��Y�dY!�ӄ�V���/rwR�ǧ-��P����T��� �V�_�l�/���r�����3�,Z���P��_g^�{�je��Kf����0p�?�<H  �!����o>DR�<�-W���0g�VѠG�EN�-�g�M��U�g���J(�ٯvg�$�es"߮���r3�͐;,�H���h�O��j�����P ��Y$�&@i��=���P*�+0�$m߿D[��ߦ��3���b�o�a�d���[�@[R��^��O��Í�cwۨ鎱Y�5f����X"N��ܔ����	��nH��O�
<V
K%�r/y�f��G`�>�r�	�U��|	bJ	����6l��}��%oQ����d�	�*;x���F�%϶�uJx�j�}?���� ��1��&{�A�ṷF-�]G��4���&fK1�a�'�a����oԊ������8J��y�I���c_E�ny)�$�����)A�
�'ff��T�����Fe*4�6����{�̤������wig�0w9sp�W�${�1�yY!���SS��0r_�ҩ^NT\��ϸ-U@� ����p}?��`���\����7��j ~�k�@cB��n��jQ���1��p��5��k����)!T�X���+����V|�;���n��v�Y��A�����j��`0���F~nы� 3T C�_E]ߒ���ec��U]!���˅�|� �̗'ĳ��#^j��٦�R�̾�'������A�g�����q��dR�[��X�`��h�H��	e�Ɏ7��z}����QЩ���q�t���-�±ݣ:��W.�n]�6�6	�CL�p����V�'�lz�b���g|5{�vEq�m��>��DP�X�ߴ\p/�����C���[��ͩ�)����ְ���B.�ն���Bb���;�iti�(��Blm���ˀ��}�z� oJ���E�}��%�
<�{J�UC��e�e �j�I���>�����(8�4�A��y5k�L��爦Ƙ]�t�[��=�rD�'ɪ���,�*ٴ3�:���G&�����ArybB�O�q	Ay��>�������6��	����";���Y�N�̡C�.R�MQ��+�։I�˪�>���w�D+����i5STR�E�<�#� �(�� ��1�R�}^Y���;"*��n[�mt��.��D���#�,��H��G���t$0��_�~@(w#�K���"K��&[U��q�GLf��o>-2Z�{�!�6�ȼ��r�G�'Maܒ�a?�L�#㾐�tsYrƢ��l��V��6����ؚ��}$~0!��,s*5��󚄎�w[1+,�I�^�'�c�P6x9�T��I��p}$�\t}{0���Z~�J����L��+�����C:���9�B@��#m�����ɽ<��u��c�Q*bCA�|��Bh�7� ��he�͚�b:'�z�&��6��o������#doZ��a�o�����%���ӠKpƏ��U֞/K鿫I�̊gm����sڽ�_Q�]&�)g ��@��ɀ����3��pHy���Nm>�I��,˘���"�o�}�*�f�,�8pI��ʷe<Gc�U�?}�����@����7�P�7�>N1�7��;=]BK��b\�J|xo�&H	BX��m�t:�e>��(O�/m�5��6xM���ÝƟ�t��r�b���
��+[*Ш�� k,���q2�[��t�����T�[ɣyHv�;8��M�wRM�o
�,���5(Ί�º�y�h��ţ���_��&�� ��j����|��;��A�5?�rMmh����g�9M�У"<W�pq���+�2��uMb���,(��������:�.����,Id5����P�s��.䀒U��MGr�|���U}��yf�[S5e$J��3��x�X���f�|^K�mH.�ͯ5nv��9+�O�#:��-E(Y'#���̹�ĩ'S?�3&�W��-�:�ޑB)GX_���C�{1����lG)�zyAeA�s��x�{��а�a{������"ZRQU�(�$ʌ�ʲ`����{���.��! ��	g�оp���DS9u��T�2�mRj�pӫ�~X*6��vC��3k�JN�LU�� oZ�L@P��#\�)�bX=�v�`�Ԙ],H3��#�·������sqX�q�6��s�i���Q�
��f�P{���+�Tl���G"+�Q��]�j�ЋD�n����F��*%�V�t����U���JU�D�5�V��uz�[2�s��_����iz~"�%:��^sf`Ú|A�8ؒӥ~�ܽL�/|qn*b���A�L�I���IQR?%.
�"ӗ �B�7 o[j��z˃:(�	!�U��y�Av_r6���K'��b��'�!��اE� �I�5����=ɥ�P�%��	u8��L^�|#��e���R�)&���N)?/�Y�Vp"^�XP�e��B���m�
�Fx��l�n�`$�ɳ�R�2P�\��x��1��ٞ�'���jͲ�����(n.�.0���!����Iq�9�1�2
je���5����n�W#�vc��#�O̙<'؛w��~�ڤT'���\Lzg� �D���>�#��N~M�#��T�ݩ�W|(�YQ�W�$�8�$�深��{�i���F.k����BP��ߓη���ߏ~P���a9nկH��H���W%���ߞ��~�k9���8�>hݘui>�p��wL���?�.C*d��KC��Iz�� ��	-�p�p3@}��we��1��wj�f����S�I�O����I����;{�����	z����T�Ýv*��V��O�s)��/,����AXi}2WA.�x���L���b�PK&����p�6EL�?�So��Y��tR�M�s?��� T�a�X�|�%�n��h�_P׵,�`��U��e�>	�>e�1�?u;1�tǁ���Gde�7� so��O(Ն�Nw}7�C��چ�h��M��`���'�=]~-�����c���__}0<c�2;)��]�ԥ��f/�ϫpׯ��-O8�4�Pɇ��B�����V��7�4�8k�����KNQ�=gMz�Z�Z.v�Ы"�9,{օ�LH(�|����ˠP	� ��Y5�M���,��V��`���Oe)�m�>@T�f����ǁ�������+���
F��iP>�^��(0J�@�"���1K������v-�wʋ���9�&�����g+Q��<Z�1K��H��tr�L�54A��f��"���cB't�f��z4����4"h
�2f�+��u����%�z�p�%aT�ךW�&���i��&���?�S2}����d�Oݸ�}]���~�S��*�|�JV�Ԏ3Wd8�1�g�_�3�5g�b��b�H$�Lb���������!%/���������q�i dã���-�j~�!M�Co���V����[-���t�r5zL3zC���R���y�:U��[�����~��f��mb���\t�$�8Fb���%����������E�����:�o �����4Xqw��H�򫄈��G߹ٰ����t�MQnp|��7C~/��Oi���J��1�KY�c�5�%mh���-�{6�� �x��B�(�?/c�?&�'-�3���"�*ʪ�>z���Y��?��3!U1�|����9.mTj�tk0�દ�i�q:��
�ߨ��*�^�񎡮0���0�Χ]���+mV�B�p��[��ꄣ�%�h_�( �?-0�_�7���_���X��ɫ`,]��ɟR,�	�܍j�����q������ ��w�Gg�p���L���K����ߌ�E�쐸�A3�<%�T�(�(��e�XZ�u��qb�RHjx��'�	�����΃�?ܒ� dW[{c3��|x{��q�A���>U�B?7:I��^���*�A��8Q>��(p���"�tHg �u����:(<�>Q����E���(�����u#����]_����5w�~9,�lg
���Sx�dY���H�S�h�M�_Ͱƹ~�:Б�x��Q��"�rO���3S#�j��L�����s"��]P%s
�[]��~��N��b�蘡Nl����ӿ�k�XFÿ�r舼]s^��4��T2ޗ|�Vi�1�sQ����|��Pn���@\r��
��I��m
�Г��^%�O���M=2T{2eȝ�pw�����o][J�<W��2ط9��LSS��۲���G�O�� ��y���w��Rr^YH