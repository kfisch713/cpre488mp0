XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��E����X������qD�:��*�����mOޗs\�{��1��#��`�����3O�\VC��S�ҁ�_�Z.+Q	�Z]_/�<�P@AO-���������z?N#d�Mj*IȎ"	����/��G����[���/eu2��Hy �,{!{8Gl	>حh��c@m\%PO�������3�v����s"9�]-<!���V�_�ҭ���,Lr�5��7�/\v�w��^�4�	0�
fͭ��ǭ�H�E����RB�ըG�/��j��\!lg�����n.c�!B�&��SNyP�; 0&��+�4]�N�ȳnO�vHE;��Ө=*�Tݒ�(%��S�C�}R÷��+��4����O(���i?�{I��/E�'�LI�����������c�5N%���T!�7����Y�-ٴd��Ck��˝��a�t�AvH���Z?j):�>OJ����ZW�>��I�B� w��5�� ���#�I���(䪍D��З�e+q�|t�"B#���+�����$��k�(����~>B+����xK���BJ)|���|&����2��������۞��i&�g*�:C��q�6�-(�ny�;V>�"Ȧ�osc��%�����$*<�Ёd���s��GZ FԵ���h-�m��@�F!씺������]b����'Z�;�"0W˺J "�Z�{U"��76v� Q~E�n�h��Ӗ�.uG��œ�nC�F򬰩c�#C~a��ck̵�[o��sXlxVHYEB    95d3    18d0�Aǆ�L��~2�B�6�H-Xf�Ca���/���pR��_�+~/�������-Ʉ����;������듘�J�%��5���X��&�6��*N��e-���d��Nl���җ$f�>�^S��t*��x�;��%
s�>��y��Oܲ��R=��TB��M��}{����xM���-�gz���Q�\��vT��Z$���[�w���⭆+��B0�X��WD2ZU����Z;C?4�G�Y	bb�Zk��Rsħ�h��맜N ��8-W���vߨ�ʯ�T�>!ږ~�!�f�[�<A"�!]sؐ1��@s(�K�(_+v4�o���N�q5q���|��y�嬌�#0��O��Ĩw#�(Yo�ﾐ�we�����>J���tEb���gE���&q���PY�A�St�Ce�`�@g�Ǟ���/��$��lV���f�e�����j{s	IBn0\29�ߢ)q��jl2ݪX+��B�`f��:6X2�P�R�O�[�>��>���6;�,pRĽ��E>�,	ֻk�SȦ�+������ �iެ��dJV!psM2��i�d���<��>բUy�'}��<urG:�r~�2�G@i�&��쨰B�I)�����=�Ƹ��A��� �g�����ƚ<��RDYr�U�d#%����V�L�:�=+�.�C�{��>Z�Jh:[�	�(��_�m�w�
�T@���A��ս���O��	�� �7�a�M��k�8��ḫ0��8�@,-]��x[�a�#�. ���~(q�mF~~d�[l�F��6��D�wU���k�j\c+yEl�����URtL�Dh���I��KG��z�,!e^S�6� ���\���*�^��Q����s�*H�kHɪ�j�p�s��nߤ3d�.���Le]c󰳍El-2��Ե�Tf�m����"\�h4R?��s�x5�������R�K�����qyI��Qck�Id�&<S݄��q����������ns�"Ky��u�0T���C
���y8�4�o�1 �u<DsJ./Lp�/B--G��ı{Ҷ���C�d+�����C�~��B?m9��|���U��e�c/�.;��z��
ɯ�G��̑�^��<F�pѾ�^\7t��f�
����(65}�&�	���Tn�2�*�U�D1_C�#��h�Y��;s�	��8�vR�ퟪ?�������b�@&��t2]gd�� y�mG���:^�,��	������3s��Q��$���c2P�"B�.1�f��>�^���x\�i�������t�T��cA�4�B�fL�Xx�&���
mQ(D�4�'#��N����Lb�8="��|5�B$��L@����>� �Wnm���]�^
:�[�v�3����E��x0�Β���;�n"nB�|v]���D0��f�Rd=d�-���Ϡ��&��FB=�k�X�v�PG���1ס�/��r�i	� ���*o�����1JP,���:Jp�J��G�Xҳb�5�X'��]��	Ι�V;�.�l�d^�2�,�C�Q��q��3A�Oa�_!�pZQ�;
M�Jowq���U�|K3����	Պѕ΢�V�9��w���eYF�:}��o�d���&à憜�~�3��&��� ���Z�"﫽�7�@H#r��2�_z��ZnZ����T�c�12�2������52���7�_�d7��W,g��6gz�=.���߫}��2x��Ü���VC����ٱ�i�S`��YAa�(y$�9���A��1�����ǣ�(�$�Ƨ14�Aj�9"�c�6�ٟK�}f��^cW��v��>;fz�1�3h���g��з��M��,���C2�XY0����'�\!<�u݊����ٛsX}�Gx=�8�_=iq1��)^�Nj�Of�"�����'l/-}���ndZ�_�$���n�h�+�}��l�ϴp�pBn����}��C��ʗ/E��˳x�Pn��ss�\�Go��d��A���ÜG��5nY��� TLʔ\��sp���̡jBJ�����$�q�z��i�a��#��2Nß��(1��l�&y��zi�z�5��2(��A��S��e_�K*5��r�.�\O��Z���Չ�x-�xH�U�!C�ΞG/���rX��ۣ P���bl8��cs��E��7�A�OG����Dڕ�?@��Hg�h�kV���8�2_�tW�o<UƠѢ-M�z0�/D��,4^X��q7����:�]+ w�⹉������h�ŰO��Le�"F�2���3�?g�d�p�Ud�0t����>�-��k�?���H!���5�^p�5L�k9��朋3n����������l#�����d	AU1	����-�ۖ~���ٚ�̓lfV����nQ÷��לRN�����eV����D��ʽH b�w��૝��a5ɵ���D{��d��{����'�m �������M�Ș��L>���a�ق��s ��fM*�$�ՙ�#��J5k����r��b�c�ZJy����a���o��7�ɨt���ww�|I�Ǳ�o
w�R7�:�i(0�s)��3	-	�W2CyEg]ၕ��l�n{���%�)2��,bk��LP�!�:�칤@����矊t��N��+NI� 3f�X@*����Yp���{����}��A㝅>�,�m9J�o>�Y1�2�D�2}���}b�'��Lݛ��oA S+��طd5���B콒]B����b��AZ�!�
��2����Й�)�h�:�Os�E���=+�3��J�E�����{@�ı�E�Cv��z3_�&�x~���K�,IS0��
U;,\�h�<���"ǎ����K�H�����h��Þc�8���4�w[��f��#+��g�*-�ܺ' `�����¡��f8^Z�}���_l�p��p�3�v��� �M�	eS�[>a��#��B2�9�\l5H�:o`I�A��"(�m`�+�NRu�_ �����ӽC� ����v��{����)P�@��R �5�Q���^v<Y,��X�f�ށ7�BP�4��� |�w�48pw���L ���9�,U�Q�M�_D�?"�=a�!5V
�����HS���xQ�[Q7)�.D-B��T:R���8*?��@�H�3M�����or"t+�r@���k�"�N��\��=���i��6��ӑ�<c����SsUE(��Ņk��b�����tP����k�z��X��u�����p|wi�3�c{��������Qg��!�d����;�tT��1*k�̊G�q��۾^7�>V����Q�a��O�Y��)�	��5�U!�{2/��c�}�Lt0*��!�3%����2�Ӂ�v�\��A�-0�1B�4"0�{T����b��-��sf��(ʯ�m�4�N:��O����01Q��e-O���V�s��������z8�?U��V�O!c,!�cm�z�L�d~�����ң���S�U2�����`Z"���>ƒ�YzB R~e1$2$+�|�������ݒ!{0jήOk��p��9�Y�c䪏�����_��%kS�5�tg�
��86t���S�6*�y��,�M%̲k��7/��r�̚��5ܿ����,.���ܡ�v�R��iS��dp���`���}Q~�������}9��@!��U�)�畺�$z�N��J�t���G�l���7F��+x�1����m�Sg�
Z|�T-�ey<tE�c격���#�?Ȋ�{�s{g'��@�aӾV��hp�����P�hￕ�X6���	�G�%�'���g�7�7���6�J��:I��
lSO�b��פq�˭���# }p]������o�����<�p��as{h�i!�Fe5�IO�X;^a
 �A��#�WgD�|�<��`Q����Ǥ��DӺ��V*�y���Eފ��P{���ڝ�mA�vcbKX��;��GCY(^��b^ea���D�}p�_�dT �,<����C�D�$k�^������2� G����Pw"����,���ju���T��{�U��$�Eoa�[4E<G �9�m���u��i�&o�)}��`����(��Wvp߻D#'�����&<tF�wr=S@��2�Rr��?�	e��}`� Q����Oa��L����A�V�6-�ʀ��1��@���.�b���ho��˅���� j/�s���uc:w���!d�U��i@�9�a��)��,o7���VM��7�Q�z.U�����ɼĜ��p�H(�ҕ5+N�IBA�̭+�P������!�$��\���h��KG��p�Q��R�S�ڸ�a����Ǥ���T'�Z�L��� {�<�E+��J���xB�Q����E�f#�û'��xQ:� ����q�-��h�O�\*�a"�w}�76R�X[����>�B?�vj�!�TY4CF⣘-�Cz�u	[�	����$�I�Hb*4����g0���@j�:�r���O�fxM�7ק���HX^}��q��|��n,�6BաD����qS�H
i�����S5"uQ��q��Lk��-v"����/����j9�?�bQ�3e� 9$�4`�ڑf�9l%A"��7��f+�f0�Ś���2�CU�c�F���Vr��tQ�=ۦ�ELnk� ��a�v����'
U��M��[�Dj�e����A�#pן���L��B�$�9�I���S�T���:#,��F~j��4a���1R����t�j蚤jCjMXIS��;kR�� �G���	6y&/�Ju���r�Vvl+�� ���7 ��+��������ݶ�sF $+ΞP�����XN�5:ޗ�c2�l����i
V�wv(i�=,��*�؅��8M�� � $]�NE
���~i���A��L���g��.��v�VC��\�
'�}��h�.v��d�*KJ
=+����a3�;\E��S�C�C �r��t[tn)A��������dv� ��E���_9v�a��w�|R�Ou)P��'��#B@����Iԋ���d�̆��%��	ײ�6~��b~D�c��B��ɪ=^�tlF6J/��Ƙkt.�׬���BW3/�0h�=4��MD���?R���e��G>�-�N�d#C�ȓׇf��Cs��i��A>Q���U��D vR�MN_���!��e�"�˦�PF����aSa��Χ�X�L��R�y|!D�����LO�u���6o���(��'9�{Go�G�;�MUkD���uӰ�!W��ZW���s��H`Sۃ�J�i�Q,b�{�������-~j��m���fm��7�Y$��r�����a��L�j$�
!�:�U�&�)���p��\�	��rGE��]�'d�`w�L�p���ʖ�����D�|�d���Ї��� ����l�u���#r8��M[#̶߱�.`�+�ߌ" ��{��GY��1l$��^(���LBw!S�kTbl�-����:�I��1�� �	�]�q�\��Xӏi_��m�P�uC��P1R�IS7�!h��|I&��&���.�,n|��F�Ʒk�t�nh�N��b�d<��De0w"���F֑�x�9Kt <f�����T��}3R�q�皑��y:5��~M�����w�1���B���+���Q��v�F�+����39��F;[͞�хa;��rD_��J�I�ܤ:�s0x��Y^����T��{��L�k`i�uڢ���'�T��mU����F��x�����Π���v`Y�"]�yƁq�.WYۂ��j�U��~�X���(��G����vt��w���>�sZCA�h"8G��)�Qb]��mg}�f폎���S�����<?
�voq�u�:p�n�XQ���6O��\�kJEP4�7�?P?) �y�m���|:����g�pX��Vx�Cd�����m��s�8:�\��{�,C�6�)Yn���M��7�2@�FZ�<�o[���e�B��>�w~S~����?���M<#^�p� �W!mL�ukÓS�dBv�!8I�	�Ri�,3��[�gB"꫐��Ҩ��c�~��i}�﵄�Xt�B��=7��~�}��pb����6ѣ���M}O�1��>����c�[�&cJ�;���w]%|{`����`@Su��.
}!�y��W%��Mz2~�i�3���A�'�fqp7\z�VV��Q���(|jZ�(?A��,$I?�CX�S	�fRJlH��q�5~�d��