XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���:������ENb�oFS�P�;-�b(<�D�0'$���C-�^�V���E`�]�ʴ�� ���}���ʫ6=7d����6�̡P�6jt܈�3µ�'Q9깁r�W5��4�d��]�2����إ�R-�FLEͻ½��*�剂�RA�KO�ыNt׾�p�*��d�B���y�Nw�N��+�D�N�f�)�$�#�ypif�͇��Yx�M���TlG��Q�ީ#�m��wԇeg
��,�Lj���-�;��v��&g��-�����9��5��+]ح��u�?+���Y�@I���W�)3jfN���7ƭ�ܨ_W	^��ݔh$)4(����f�	�a�h��|�訧�'̻q>�X�0������� �"3�>֦�j���D}G��{�w��0{�T��hNY�DaF޵
��l���&�����$����r�>���Y��H
��i���-��,�2��\���ʯVL�Ȗ]\\{d�a�)+wj�Ƹ�c��s�� �Dϳh+��{8ŭ)�%���W�l�uY���M ��b1�<���_.��Cƴ�W��N��V�噮�C_M٦�� |�b����_p�i������t�9�W(R��_�7l��c�� 9?��-�aZ��ŗJ�6�A�U�E<뾶c�1=H���}���}�R���S�\?��EٛΪE�L��&��Y���@C���R��;!�u����2lJQP1��	�}I��'�?��>ś���ʱ�<x5��ǧ��3�XlxVHYEB    a037    1fe0�1ns��Cx�w�����1���(�M;'�4���C�O�a40)�@��&��}A��7Y�b�AQ��|�nK��S��r"!ܺu�%��x
;�!
��i�Q�O�3/مVM6l�ơ2p�j۶��<��qw~����?u�6�bٍ�tv#ȟ�u�#q�7- h�E�M�����:�J�>��!R�%�&����������FI>B�&�Q�PtȎtxG(an�#��̦��ڭ���C71Ŗ�[:%��2MU,{C�d@�K<�[��g; �D_-�W9�����x���Qsq3�J�	+�  `�؀��Q�a%�/ ���Vߦ��,�dt���a{��
_��� 'u.g�]�W���9�^��_cƝ���<'�|��i@��@�l���ڣy|X�X��wb<˅TFB!S��)*�5�{��N����x���	%b�X�b��n��qb	F���7�6r�,�?�"����E�΀Jet�O ��SbУyH���Nn�kmi �bxur�W�wS�"�Nz��"��.Q�+�	�q����O��1�Wc��j�)�H��V���݂ZF�0 V�U���Dbi�g�T�h|LTnG��1PT�������mIx9�C�"��4�ŌA��h���<��F\��������aj���H�5n�~��.��(���������N���N�K0��Jo�|ZGG�[�N��R'�>\���:�AkD�/�{��*�;`�O2^�L��׽l�b�u�?�`1�ν�^χ�Bm31h�z��*v�G��l����vh���ه-���?�a�A��L���9�Ͼ���%��C����������gn�����'I1+9���s5�.�E��V�H|�ι�ꀅ�
#�5��JO8t �U�̼��,�Ԣ�(k��̚��AY9�B`Bo;`o!�{y�u��7��Љ�;$��g_9s\�zvA�j���U\IOYG�Z4��E�]25|��"j|�����'�J_�N
R^���>-[S�Ѻ3%�9t�"���%M.MF_���f�2�)�fɰ������{�CP�:֞B!�CN܉��Al0��s�qY��Ev�s�@8v�{��Og-���K�{��UW�H���H�	�"��]�d�ǉ.jɯ�_�����A#�OD���9�+�[�������{jGB�j��t\qmD���|&�J��ɵ�"�&���P�x�^.SC�$>+��������Al�0�O������������Z���k���a,L*��8	ae�si5	$U���Q�N'Q�.'��סv��d��X#RUG�{/�����ۇ�T4:���zJ������4ߍz=y���xHuX���
�����̯�l���w���/26�i#v]pm�����r�����������I��s3b�$Z��:i1�ٳ��4�̺ș�./|���Gr^<���<�F
���Y/L��"���E�%&�K��g&�~޹�"�fٙrv� �q��H�M�x��Kf3���Ҝ��V���Z^I�v�n�o�Q��_\R:�A��J&�~���0�:X�b�b����]Y`�y�_�;#˂�܊�ih	�F������|��&�R� �X��Q6�^_����~r~�� ��O,$]�~k��j�Č `j7ʾ�&z��2�0����a{/텟J�\�O�y�/*_VGA?^ CT;�"���h��p����T�����U����m!��U]���/U��BO/�
v�����e/���ݛ�$�2kx)m$�����0ۤ�b��$]"m��	^}"���R�u������S���\@������{�����^�*{bД��ݦ�����H�
.�܇�Դك��c_$��m�(U?��j)@W�Mf�H��z�{��͕|�&g:'��qT�A���8?_r��Dڴ%��ƺi:�_~E֋�����2�/����q�d��KL��گ]w<Y��e}���ɽE}� �Iy��	����<��o��`��WR�eg�1 ��W��x���?z2jm`ϐ�����w��s<,ht�snMM�������y1�J���nR���k֔�"�����Ɔ�d+���%s[٪�n�(�-����i`��}Ӑ �	��+؊������7���l�4�\���e��t�Q����yHOP�<��G�,܅�����Ǘ�zK�\1p�'��p�V׹�(Z����;������Q��)��}0k�sTj5����KH�&�.�AKM@eN��H%���ӹ�(V�i�"~�Ģ����es�Re&c�D�х��I�Z�E���L���b��������"׫�K7X底b������ҥ��7s���;?�0*h ,�U��F��;��bt�Jy$��]�*�������M-!�R�d��	^��v�s��Ln U6����Y������̛8�yI�G]��9=~Z���*�E��ѐ�F�aNՋ_�|�r�E���>����K��^z��ϮG=N���p$���$рK�B���R9�`=?�`��i'�6(�Nl�5����C#�U �Y&nB�_��{���r�gX3�������@E7��3�kq���(��\���A�iz�w{�m�A�Wĳx�<ߴC�#p-8�t[q��D���	s0� �o��iK�К�-�G��H§������WEZdFSZ� w��T�BZ�)����Bڛ�RG�	�cU�g�-�w�"�ǐ3n�jvu[9�g�.fd����FEZx~m����2ߍ^;xo
c	�>�%�å�����i�lz�)>0�]sO�C 6�%E;Cf2��+�U��b��hz�7s� 79��G;�>0�H[�μ��5�8y}*�{�ط��K$�MD�^C�#�Q��X�W�_��`��������:d�$i�.�ȇ�T��%yܚB�7%�R��C���B�	���48���ۀ2U��f���s����P�����Ҫ�x�h*[���$;jPkon�^H�Яe��K�'G�bM�Ǽ�yz; 1���8�=Ԍ������h��/S%��Ю�<
jKW(1/^�(�����>D�v�+��hL�YX/����@�!*\g �F��)��SlB2���/Y��#����}�|����ӹ0�'/jy��8�1�ޟ�-܀[�ަ���U��87�d�;�'kv�OW�A�E�8��"����[�����O�5M�#��.�AD�ξ3R��.N�.�k��X��)����w��RALQO��e�ޛ*E-�ʜ�v�]��C�/<��
�੬!�� ��܋`p�]�p�'�����핃?n�P�߽]tK0���S�eoL�j��c�6C�_�;u�.��=�,�8�Fu�@����/�EW_]6ƽnO���no3�C��g+S���묧Uɜ��Ӯ��wߺ`�v�$��9��?kgb�B�'Oiҏ�-�27�i��85j��+�N��r]�c������N�����P�����~h�ؿ*	�1�E�c��؄ L�}�s0%�?���Nq9_#�7S��/`\�E{����%��K!�?�� �f�������Щ�fGJ>ʥ����_(Ur��[�c����9�����7�/\����g�6��O���1f��c@v�z T]��e֡���Ԣ	2�����u�P#?��Pc�0s�M9����\���X�l_ݜ�~f% ����ee��:��Kff��@eY�s~�0��
��t@�ѣ��*�D'Q�HK�vР�[���~E�3՘8p��;�}���,�@�_*���ٺ���iW��Sl���E����+��͸����t$ ��85;q�8͸$�(n[v	F`�	*;s�n���=h��z3e����Acgiv�~��'�ZCC~�Sb�i:3b�!$q�^�kNW�L��녻B��F���|f{C�\}��륵>��i{s�$�"�8u�z	��*N��w,]eP��>�����R޷�c�9�I! �����="WE��vΓF<��44���J���=�Z�˫�ǲ��(�"���h@����(,�kU<�u�Ԍ�b�4����j)�I����;V���lLhܞ>;�wW̿�Z-:�I:��#"]O,�D�� (�*2?}�^E`U���e�}JCs7T�-�$I@�[m z��Ď,U�a5Å�灒wCW�|���w��ڹ��"u��K>#�{�wJ㣤%� M}�_h����/�duz5w}�����;+�Q��*�_�,�sv�n��c�أ�=�g R�^k�����JGFUW��2�x��EK�����t���%�hW��s���T�1fիJ�E�X�I��~�)\�=��'�Vy��v-����?�;6i��X~���x��H_��_P#�_uR����Xͅ�$,�$[���M�sh�>�RlyC�������:��(�0l���8˷.�A�^H<m�E!�L��q]SC�ꥍ	n�b�B<�o��)7�{Y>���c �o�p���b�sc��i�2��]r:��	���݁�vts�`�EVNibpg&<|t�z<��=����]�%�>5��mK��(-���h��{'s��\�\°S��qQ��w�0��y�@j�
�6e�Ia�{䑨�hg!=Ҩ��J���Cd,K��ә������S~��Ba%�hH��A�v��:&o(x'�mCjyٵ�F� �1�ө7�w³�J��6z�r���`m����v'��tхꔄ�g�	J��7���z��fO�}�$�o�pj�ÊF;�:Cp��������Lx���ԑsp8K g��ؼ�0�!�|���Nq���R�^���������Q�m{])��W��tDۛ�h����p�����$.��
��_I&Q�Ϟ���������g�l'բ5R�C�a1�`#&�SOq�Q��ٷ��-�-!SUp�����iځ�K�U�`�.��L�w��+e���?�wv�K�^6���)K2ꆡ�d��A�A�<��#�	���&���š >גl�e2���A��/�&� ���y,�lX��7éD�0�ԍ��� Ž��G)�C��Z_,p���nq�'}�\3��)��c����BwT
)	�D�m�`�s<%!)�SC�G�-�>��'�s��;݂�v��^2���ʹ���I$l�ùt&��uK]o .�e����DQ-��K�#C���̑��CË�G�r��=�-��E(���7t��M���[��˭���K�֣V�#����!�>��FH���7`&�ߢ��!tc����F��0���%��cK֧��w�z99A����kv��ku��U����ٔ�X�I�˾���#��3OE����_+u���3�z!u��q�z0��3��"���u��wV�ub���ᝲ�C^�(V�f�`��'�k
�2Y�O.r��K����3C���}(�7Pv����邫��O�G�=G��Ɗ��g�ۏ-C����L���)2��5Of�EPP�a-{�{��*�r�SP�|ȓ���u���������#k�!�q=Om+_F�:e��@6�f=��g�������}��"۸Q����Jؐt㊠T��������2Z�?�h&��{�(��[�`��؏�*4\��\e1vI�Ԃ_٭�?"�P�<vΟSmQ���>Ex8�2*�J�J`D���aڢi�V׋�/�Ȋ�m��N�.�͜Lվc�N�_����L�����tB�E�*��݄� Xl�g�R���r��@&� y��xR]�*��\���b$%-B��� t[m�+� >.�IOĨQ�d����]���`�ܲ��2�9�I�ʶD�\��m�|-1�ep{ռƢ�Q��DC�csKJy�@���&Ĕv���b��x`� Y`LSl=����d��H������>`���z�*������݌�.�Gul_�SӁ E����/ƃsKR��1ԉ��(��Q�zZï"�!eF։2�zc�F��HW"'R�X>[�O`Z�_.
��$Fګ�6�(�XCa����2W;Vz�^�*C�OA����z`��x����`�Rp��&V�!%�U�T���}ӥǒ�`gP�a|����<m��-������[��o7'6/�`��|�c\<��v��������>��Ԃ��������=��ҞIh�.v��~5H�z��h��
���٢��!�R�|�r�ei���N������2���|���Eaeh>�y�����ZO�Z@�J���YCىX]ޣ�SR��S ��Ui8��X���Ѩ6_?�O�DCh�44P֋�#�����I6O�WG|�s�c��3#�*ڦ+�6�R�h�`LU�6���Tls}��:�U#��#�j���V���c���DC�
��C�ay�X���%�H�յF�����w-p�_ ���T�-dT�����v=��!��C���y�B��P�װ��h�'�wObjs�VjNa�ymx��[��@ӆa�c�}����y��5�zf���Gl��ɷĥ��<-1$���n�C��Aj��V|��6�z��QI���=Y��~��R`\�C�.��E��@�`�I))R`R^�BJ��^_���d_��GnC)qǷ� S�w':w����M,���MJ��9���eg���Ɏl��I�٥3L�T��5$dVQ�m���z� čJ�s.��4�����aϠ5���� wM:�-�/r ?<�gh��='�	��\��H ��h`F�aW˞J�y��Mb��8[|�/v��^�Pqy:}��� �ȧ�pa�tĪ�m�Mf]A�0\
ry1�F�ٌ?���8%I��Vﴢp��Y=�yYu,����ci��~4��y#�]���{��ȋ7��E%����g��$�"����_r��l���֤���}�:u���ݻ6�k�0��~(�fC�`�ɇ7�0�(��.q~D^]��w��nby�rop`;���Jv�����qT���n./�Bm�OO�:��o�ۖ=�u:�E�� �]͹�}�.��y�t*p�?a|�[j6�<.'㜿.�J\n;K�2�Of%a�0��SG"AIڟ�)�F@��U�r�,���k�I���+�v���r��st�cxn7�K��ۉwJ��x�O`u�b����B�I˷d��jɰ(����$�xt�
��j�����w�6�U9��u�'���A�lB̿�b����Er���(׏������Uc>��̶�ښ[9�b�@"��^dF;B�&��,Ľ�LAo(7E7;{���tw�@�EЍ�7_�r7�lB�/��ƫ���W�O.e���D�&y���������\g z�l������X!E<���yt��Y؉>gf�4�M�����{�5o�V�tIy68z�v��=Ic���X_��:���]Q��)��X1���PRij3wq�н]����~Lf�H��/�'���u�|*.҉��_�.��w	M��7�A`p�]����h�F��}�k��#TQ�Yt���y] iz�8��̸������q�Q��]�TJ�����\s��.����=��?+�2N\��߇�p{�����]��{�'�S�P�}ϣf6��e'eR�<�����%i(�F��(q��%��gw�MK�}nu�A�,���+�-Gz��78&+d���3r�o2��;x�$�Uy�J�"i��'����M�v���2=m�l�v�z���M�ݝ(�_�rl�w?�6OW�4$��{�B� �r�ڜ�����&�V�#���#?SU1�`�m�Ky8��Ȅf#�.Y}�O�-N���S�kRI��<�f�]���36H�9���fZ2���aY9�V_Hb%��h�\�06��'~tN�$ڲ^����S�^�3�v��?��U'�$�V���3�yA�[�g^0�,Z�0(���R��`����qnrZ�Ytl>|�s4Yufq�2�z���#|(�_:Q�-e�h}����2���PCn�"y�"&���ñh�<��\Z�C�k�&��<��ji���B�����Ľg�0���N,f�ZJZ,_�0�ɳ"����+��ʜ���� ?��_tun���y2�q	 �1�H�?r��U�
 �ɠ>��z�A�]�Զ�,�