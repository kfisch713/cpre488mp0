XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>hv�r�"�>m�TDU�# � ,���潹��O��xr%�|�!ɡ_u�R�BZ��r��&�M��_�Y���¾:6�.��ˣ�[E���H?��uu&T���bd�!��p8�$�<>�]���;���_�T�Qe�K�	��&>�z��h�n�ly�@ ƚd�`��6P�����\N�+�&U�̦�+�`	�v�$t�N9Ө��@E�9[��9Џ��޸�x�E<��j���)����o	ݔ�$\¼�.bg�s3:?6)K�@�y�oZ�7yG�� �*�`����ME�)���R��|{���w�_�;|�����&��(��U*	7�^-fo�ǻ�B#�|��{b���·V���o!=��q��c�9y�-��j�+�.*͝	B�u�r=Х��[�4��AK��$�m�K���x����5��X�a�JeE�$�b�+�뢮m7ڝ�zr��[7�B�<L��T�1�J;��ښ8�W��8�v��د{�j��[�D�W�JG���m���݅"16<����a#۾�/T�74����C�ˇyVW�"�!^ś�b�:rW�"(1�d|?
N��t���7�Q����\]F��4���g`�3_V�h���y!	� }E��Ä��y"b�*[97?�9zWĕ������1�f���\��n��c	HG�ao�O��p��e?T}}�oRv>>M�Q�ⰺ_�ܴ����0���*Tł�Wc�����b"k���H�6eS;�OA&g�M��XlxVHYEB     f6d     6f0b��Z
ϲYb|UX�G4��-�\���
�U�Ȫ�V��?�R���75ﵺOu9��ꪕN�_j%{ڬ�1�o�Z�V_�km:�n!�,�Bxߐd��z�&k�tW��'8	n��{����`�3����Fe7ȡP���Q������NZD�│,ɝ���xeD8��<nN��D����R?~���y
@��2�jOp�]���t�t��m�m��PU��K��d���nYh����>ร/^��lp�p� ��d���m��~����6)�J����c`L����9l��������O�� ԧ��1L�^74I�0��0iT� 6V~�)iG�Ϳs��C��G��?�q�S��|��$�A��~��K���C� ��0ޔ��k��}�;D�J�}qĪ�ӊ�˩�p���T�ȎW��t�N)Z*�7�z�k�T��� ���w���k���Pf���Bŏ��� �+��$臨�Z�ͧ�����k��:N��z�:��nZ潉.�0���������/G;�z[:)ע%���FL��d��i)�Z��R�:�r�dN���V����T{~�h�v��J�`?߁	u�H�F[�M󾎲~P4j#���J��ܨ�.+ǖ� |<f(~և��@���Ά(�,`�G@�]��4��}��v��(�nP^�\3�Gr��+�N�MF�PvT���r��w�3w?�0qo�W��S֛cL���QPg2��Ox�v����&�ݨ���;���V�(��q\W���Fu����:[4��v63u�/�]�y��
I9n���Zre���J���r5�/��(�YR���ͱ�C�:<۲=�I}���\p[-#C��@�tZ?�X��,�V��B��ށ�cDܭt���jyi��Hs�@"D��3�a���!P H��|y֟L�)�Ap��w>�u�,���� ��:tV�{�Ε[fB3�ҝ�M��rM�g�9�Ҩ�P?>��k3%�+;��ﷆ����3r�#of:�v��]�Q��q8���:�nP���(oW�j]�
C�{W�V6�#�N�_��l
ueC�sYJ �@q��~���^w@�P�/��(�9�y�a]���~.f�F�r�J��l�`�5����:3N�0�w|�����Hl�)D�և�wW�c�׉LL�*�ܓ��|8� �׿rX ����v(gԲ"��/�
r��1c�~��G%�~�sN��J$���v�Ɩ[�mi:E�|����"r5e(/���������qVN���ta����KE�u����9��5�����s�8?$V��	.�����ĕ
zd2��n�\r6 ����uֺ���%�u�} 鷀6�^��n���=�����(L:�i���h����er)�̲*�in;�K�rؗ�~w뫼��s�}-�������wgj�%��݈<ix1ƶ��E�2��e�+��]n��gC���PNh�=X�L�3FӢ��ReDM��R��y��QM'N�mN���������`#����[vM�����0*�;r!�,��b���Z��E{��F�o�xh7�"��&w}���N�'j��o�B�EQ:p��?�����X�2�D�r�v�E�඄���5/*|�&�'99���C�a�Gȃ߃�-�?e�=P�p�0�֍K���!� z
z��d �⇜2\:��Qr�8�0`�m�{?G!4v��2kE��ݡ��Hz� ����� t�Uq��$�]"n�c'v����IE��.ݵ9L݋p0�IX|�����l