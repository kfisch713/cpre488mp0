XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��	`&�
8?�M^����?��?�5���k,����R��?'Xx��j�q�.Hj	f�=�I
��[:鸒����/l�qo"�������&����F$h�{Q{g;�F�� ��>om4P֗�'��������=��)���j�>��^���О�vd'P�<R& !� '��X�� �m�VM8���v֤���?�g�a?���:��It@t ���6�ɘ�nCMvbs��;��x�g�^���^sU9�x/3L�>%*��C�!c���V��i��@�⠂�p.]/D�d<����A�'�A�"s2�kM!A�(�4}���`���BpgJ��ܜ��-p���p��]���sc��SO�\j���u��{��F�>..�c Ǿ�}C�n���9���=��G�0��zq�E|VdqY��t<��C4��}�i���h5��P�4��B�V�7.�Z���vU+���x��~����U�c�F�H�]��3B�Θ|8�HZ� s����^�
(��Dnx*_*�eON�wx=s!E����h�k Usġ_+�J`F&R�RFԧUX���J�ٮh�t�t��q��t���S��{N$�D��&�0�`@��{��զI9հDh�0�ȸ���o�t��gT=,"{��G) NC�"�$�T�i;r�8�FP!�G�m)��G{b�h��\֛)��4��+�]|�2�o��Ī�=W�:UN�`�P&�$C��S�!�T�l�iE��#���r�����l� `0P�XlxVHYEB    95d3    18d08ˡ�1)H�ь���ׄf�w�E*U�Å�Q�y�Z� ��f�闲�%j1�G-6=W�+V۲��:V��\6ֹ�O����;M��o(."w1�_��^�9��/	`�^if���!�I�Е���җ��+�OG��s4e���A�^-�Z�F����6������ͨ
W[�� �P2��*����L��?</H�[sys��A�k���2�<�'������i@W�N�k����5C6��t���'���72��!�����Ӵ��4��C:ïQ�[��l2���?��0x�t��*�ض�,==%�	�@a�YË�r���]��(K��A�QB���B�Ɗ��;e�B`Tw{�cNz~,/~��J/�g�a�k���BI�%J��WU~�³D��}*&��c���B\�I�=PL���G��꺄��#f6������J���E{�j.�	×tq}h�Wʤh�}H�sO��~�A�x���`)?S˸\Z���Ф�/=hkd�E�`�� �Ł�]� D�6ǐ�����7)����[Xu�EF��mv�דHUQ��E���Y#X��e�h�o>�r*��FƠ[��+�bN~5���y˽��L�.�-ss�c� ���I~�[��/y�+T� Zp��\�.��dC6:è���m�1�!}ik��lѢ��M�Y!t��1�O�+�P�uH&e)��r�U	;��r�Ns��8J�n��(�3}��Q�GX��B��
��tn?��e�$-#��moY����\<E�d��l�.+K�Z��cw���C�����c���M��e�5�S: /��7��@w����`��@IӟDS��_�T��=$�6��Ġ�#=0�c�/�q���>c>����OA��P6�6.}1�	�x��0�d���ϸ��~�i_�`x_30��b���q�L�bH���M6=1�eCfE�\4�fL�"�Ӹ}���L���\hn�e��h+����mɋ��[EC�n�P�m�s��hz�_Ǒ�/��зC�ַ&'��,^޿Ԥ�A��I���u�t(�`�/� �c"=H���51�%%M�¬M|�����m�L�=xL�;�ְ���d�*ZG\��J���4��FʔMɍ�E��J��סq�7aV�AN	@�����%����YW�d=�W�g�4z�la����2}ѫH���Gձ��I4�O�v$X'���Q�6���up�Ci�j�Ύ5�N��-��U/M�Nk�9A��o�����)����FY2��M>7֧�c�x�*�RnCF�`�K{����V~h�l	�/��C-����kj�_�h&�L��a��l���c&���$5�I(2h��C�l\��g]9�a䎯��;m�UM�&�w�o�g{j�k��/�lU�f���-�&��m��������7;0�h�+�5y;�Ֆ���#���,�>���Ѯױg��e9�+-�.���V�.�G�E�ub�L��wȺ�Wj�9+����K��0?6A��t �;�H̦(#_�Xy����ҳ�g�S��0ܟ=��@����6}Muc(%�-��e���!C�񏘵7oh�eA���8��6v�(�W�����I�m+�f��D��Q7��_�R��"@od2����$��N�LQ�
��J#ڊg��-��txY8�k-��k�-�WȔ-wENH���.�;;�Ͻ|�:)��%��+d�#fD���S��,`�}D�"2���3ɶ)Z�Dmr�&G�.�Q��\�E[�� NnP��k�u�����FpA��#M���y�z�jWk�2��*�LR�������f\g���E�F�^e���!l���Sj�:�EI'v��#�u��,��?1�3)������]Ĭ�*��u�BƋj���.�� @�f9�Ǉ�^�*��i�=���N�"�SZ���ݒ�v�Xؤ�)9Kz����s��`H�ɽ?�[���% .g`{?��lz!f�h/�WۿS��
E�������"t�y��bI�jA�5�����gǧ�u�b��d������G�6I�����x^���=��q�@�&�9��:��[��ڝ+��6V�С����0�T�-V@N�bJ��@��2�5sγ�|����M�z��+�:��͘�J���V���nF|�P�ݑ�� �ObHx�T��h����ސ"��x�j���`64���}�wk�X�H�{�/���3j�������3D8�~`,��E @�+�䁕/i^����sR1�����xS�Y���3��D�<nW�F��MK�Xy��c��D0Tu z[=�6w���%�v���ҋ�l3pg�k��w�`�qD6��>ĭ>D���f$_�4�^�X���mu`$�z1b@S�8>�1J)�i�+�Ԏ���HTd>��v�ߑ>2Ry��4����RƢ��V��������GRO�|��v�(��1���\��x(hCm{j����S���T�Xŀ�6��2h�Dh��է/w{"�IK ��KK@ޣ۬t�P̓�������h|���֠�a����;|���)�UJ��$��E�َ���ˊK�k&��p>��~��`��!X�J;�D�5��tz $�X߹)ŏ�����������WD�֗h`{f��Ū�\Zn�ԋ��I5-Vg�dsZ]��P�;�'=X|A�QA��4r�*���[`���+�2�ŏ>�"F�uRu<��_n�o�i���v�)�������\�iA��f=ƶM&���%���e�p��h������ΒF�bˀ�?Fy�kH/i&���[����_�G�1-,���:��,�{Ƴ��Q꼊���n+�s��DK���HR�#�\��Nz<f	~mjW"�a�V%�Ӝ�iX���Y?�
d'P��4S�u����?�9V%�vc�L�n��?|U�D���c�tv� .�N�j0�¨�4I�HhJ��e@)�� 44��cf@�CH8�W��nE���NH�5KQ*�6�4v��b�y�Ǡ����%��#�$,7�� | �u-$NEg1e�`�����ow�b��dZ���|HP��Kll�&� �0�J��Gϩ�4/)�1�ඥg������	{s�O*"k�N>{VU�c'��hN�I�>J��A�(�ڤ��Ixb�t�T�%ϱҡ	*6�g���Y�J"K�N���rT{�Z�V�ރ��{9;�#����D��Yۉ�Ћ���4�� ��m�d�R���K�g��S�1���N��9�khH�	�"e{�=ԝ@?@ �� ��WI�8I�U'!��z�^�$��A=z}i�f��>�:�73Yէ�+�%��vb;9���b�y"ֽ�S���^`Y��UJ�չ�`*�&�nT��G1ayc�M�[��k���o��?a,�X�6[; �ǵ�OM30�п�K�kq�E��O�[?.��U�SF��
q�َC�5�:QOm�x����2;:��H��3�����p���W��������=jۯ��Q�K��EPd��(�bB.[�ʁ&O��.�
���~���o������<��2KCs�Ν?��%����/����gA;/w���(��Va��Q�YYN���G�\Q7��Z�@��v�3�+o ��Ã"��������@�ʯ>e|I����^C[�瀔y���Z��z �ֈŧ��+Xw�}Noˁ�/Si�Ũ���$���#r��E[��dШ#��wݾ/�1?t����w�gb9H(��h���$H
����Yo��X�&��u�3��^���l�d�u��C��jc��g�"̡婴1���&�K.>Nʼ��OIj-Id�ꪌ�5���\x3fǈ~��砠Y���8��u��02�ߚ�i���U%�_�X�P�H��>Τ���w��Vx�O�gSMxN�R��ؖa:>����d=(��v@�ғ5�3�.�R�qu�������p��������`��]%mw��6���&~ϡ<}T�c�af�[_�����~���Q)� R ��>���+
��֯�V���v;�v(��AtU�����9���%���h�a/�9ҷ�Q��z�W���Zn�ǒ����ܤ�3��E�x6
.ªȜz���
�Rĝ�{cK{��\FUM,���ȡ���y[�m��۸���/�h�nM0��~e�+����~�����@��\�ZQ萩�^t\���0#.
����N6��T� /���:6�dڈ�{���*��so�w�N}�A��P��=��8�v,���]�{0�`�B�3AƂݪ�}�)%Y��%<�S�w�-�Zۣ1�2�Y�®�H�����(���e�;�j��jPeok���ϾòE�RP�g�c}�u����rl�i�œ�$>g,��0�ϡ7�~֓�P(���8�P����51�أH:��g��k��f~"��*��)��T�����xNFL,G٣o}�A��qW$h��6d����ԈV���x$�)���G����	b�Ӄ�Sq1�hgW���|�ZV�&���/�=������L���^ca5�
�:��ƐN��\��� 2��זR��	f���wwDFH�.��6���~��	��W�����
OŅ6#�w	E���ٯ���`�1 ̔η�l�o����d�IR�|+?���
H@g���ٟ��>��'�<Y��n&P>��"T�I�Z^�;�[(�C�o��q�\�R��F��#��V) �H���Л�,��;z3&?7۪Kԛ%��ٟ�:g��ʳ�U)�r��~��������*g]�\����]j�̨��2R�k"�í��%�9��ծ�|���ϝ��Ͱ�K�f��C�C��R#���MY��d�{�)|�A�B�� �Z�B@��U¹y��1Ҏ/�a�H�w�N�\>c�� Pma��2��P7���n ��R��
�� Kt���:�%��9|���Hf����{��i��ǚg�Rk�cN��@�xr�!N�Wӳd�=�?k}iM0,��5�֭�Fw� ?�g
󝢫�$�c�'�ZYۍ"J����/��Ng�':�3w�,k�:�t~��k�RC�%0ܷ�!�=��>-�a[ �~k���[tu��ǼiDUC��ץGߛF�5)�^����\aS�A'y��'���/WJ u�Xkƾ1�81�ӱ�;#�β��NT1�-ո�-ʊ�E������hgZ��Ot2��3D�(p?��;+��=�{!꫸����&�+z@6�>�����にc�K��0O�{��30�[��ǶHٜ"��#�Y���'ͪ�(�L&˔���r���z==)�j\�,��3-��!C����I���Ly�g�/I��:�P4����&�>c/:�R�4�_� 1b��Ӡ�fHAT���B�]�	p�v����+�H��2�@d�Ɖ	b&V�S�X��7\���I�ʬ.���Y�3��T�ҫ!�i؁�8y��OV&7�R;9,w07���4ױ�+�&"�UQF�,��`y��]�DB¢�O쉀���(����V]:�"**�0H;$�DH��J6{�.ψ��T1T�o�Vh3���ǗJ����Z��V	��{(�ɉ{���+�m�<�A+�z��e.f�g�T"f��?��|��S��K��FA�� D���^zOv��K��&0��4�����EJƩ�4j}����������?v����8��t���C���ְ����mq��:�J��ʜ61�č+B^�Z*�~��ݿ=5&%��>� �	8�J#����cf��eLC��U��q�2��9($�c%��_��nܛѽ�qD���S/�Ac���}	�M�e� �e�+iCi� ����6���V'YD�J������I�X�u�w�0�+����\�9[Z����B�s�L��sQ~}<w(y"���zBF�Q ֌*��M�&i� �)��;8�����S9*ף��F7���/PW%�"���=�G�\��?���`�|�D;�9QUJ�w��q�7R̛ZmP��xC�;�lN��)gn
��a�GP�ln!���V;�1|�mXzt��Q����7Fm�\����W\� �՚{4�@�ҌQ�����������y̛5)���A`; .A���mJ@�-�ME�Գ!�Zv�nC#G�^Zw9;%�W����0B5�8M��(Ȑ����y�-w����0���O���T|���-+�e6�XD�Y�@�+��h^�ֳ����D>3����i��b&^�P8���7Psm?�D��sɬKc��&&L��s��3#����P��E@S���m�v�����WȨ,22@R�}]j87u�ׅb��2��.3��c,�2����x	���^���s��.i���w����NL�u