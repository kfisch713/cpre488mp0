XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0r��c��p�^��C�=\��+�4z�`�f�T g.h�z�o���G)d���'��a�������;r3�����QEΝ���,�q�cr�j�"�|�"q:�&�9	�z�|����"*fplcYb9�@����RӨ΂�Ye��$�t�D�$貗�$^R3���>���_��^@N\�vJ�V|�?y�2�.��������Onb?��F��UJ�TU2���� �"�>����%���6��r�|\d�̷j�K��p���Wn�g��EY���sA�-���W���R�pX����Em	*��gJ�r,z"N�]�ٕ�Ǒ�硽4��QrK�X���	��Y��4���B�F�3*7�R����	E�o�߅�xeDC���.���.K=�7���475͹�������2��Pqd��6F�,\C��� ��&�&d!� ��.�땒H%]��4���B���-TQ��fG6�@ێ|���b;�%Hɴ~e%�n���;���<�̻<`�2�c�T�K�@���$MR�"�?�A��@����+οT�\Y���3oGJ<db��$(>VG�������]vg�H䷒�֫�<:Iٔ?%��II�מZ!x���G'�k<�"ν�{�\� �e���`N�8�����!���k��31}��7��T����5(Of��k=jC,��jC��5cbܖ�ަ099��XN�I�y(SؑK�z<5��o� ���T�qp���So�����J��Z �����Ѥ�XlxVHYEB    dd8f    2160���ُ��ʰ(����h�J�D'-@T�1�P�jF�]{����Er�V
��#Q�0b*Cj�:���p���˿��L��yA	�;��n��LPG���U�+�����O��\3�S6�g4Sy��^�<*�p���aR���u\��պ�Ό�b�^�2>e|<��	�����N���]�V`�k1h\�ʊ��3w۟�f�N�C��X�}��s��|�^�-U���&l*�toR�ŕ�j(�8>v�Z��Ty����� ���
l͜��Aͧ_%K�R	� �A5䂦��V��n�B0f����%J2x%/�u#F
]��|Ƶ�z)���t	�V|��ږ@y�J]�p�>�w�EZo�m����_%у��~3"�xԍC����t��C�����	�P��'G�M�Z�J (������JUϧ?>g����V�8Uaj{
Y�گ3w�C�q�]��T��3���"G�L��tF-�Ik�Si��f���V����W�+�Y��j̡B=ȔM
��ı�@��';v��:Thw=�{,V1��B�kw}_-����F=_y��H����Bя��O���K����)�i�H�bK\`?��m�>��ˑY/}���?���w��1���8m�����#�4���X��c�t���[{ԟ�|���ӣ)��s9���x�쓉b/^Sk�w���+�����J��7�i@���-��G���k��>�\Z(�e��(a�(���Q{��͎(yCA������_��X�A�&X��&��Ё�����C�G���[}�gu49���V�ִh�1�������>4>������&nArVj����-<o��/���兪��z&&J�F�g�k�>
�?;�O�2�Ѓ���Q���x#��g�G��h��z͇�~U�`�fX����I���<ף�tM=Զ�˿�0
���i2 7@��@��D�AW"����Dch{��7,̰��c�1w}�{�[�D.g)�8�����'�G/hvIs|����j�vm3ǔ�O��֣�K��4]���.�)|�m׶��֤F�"��]���$o[��=�ΔD3��Ols�ع���C!ŧ
ñ�ͫ�͞'����[���# ��^��B_J�.��CJU�{}`U�j�-�ԛS�x+��aK��|~C�r�f�lJ���$���[���C�TT]B�f}��h:��H:��@F�1��U�2A�^�E����%���v�{����&E��9r�שi������U*kz�\mo0:���X��ok���[�(2�&6M��d�:6�2>7ۛ��j:�,�w�ȏ�bC6B��K�4Pq6����]�8M�*Ol᡹��Dh n�<��V����{��&��W���z����su�w#�A14��$�&<\U�&����W%�Ϭ
�a,4}w:�yۚ�xO����=��C(�jQ�ru���U������P��DMS^���huDç��i���MJl��RQ��p;��9�a��$aƔ���zeW�<���r"�j�NaF�G�h�d�݀�3%�̰���Ty ����5e)y��+Α\�4�I5�3� �.��3ז) ��{����I�����$D�YP&��Q�H[J5��$���G��Xq'=L�}���M7��M�����h@��j��JK>��H���s����dz2EҨ�B8���	.f�f3�߯���R9��E`�Μ9"�rTf�)�e�ƫI��1���}�H���; C�Z����0�-��ı���~�/�Е�,gY�Y��_���+=�Qi���Fu_�ޝ�J���j>�wvtU����
�qk�����]%}/���O�j�.郄�̌,�_��ܟ��G���)K�ErB�+̆��b�d��t�EK:zi~���i�ڪ)����:IX4M��O�\DH-��|����M�e���������Ƈ%��"w��_	��́��՟�����"p�Q�nۻmj߼W��չ/�C�gd��Z|��� �n�o�=
#�Ϳ��~��r7AA�V>xCU�*O�uw6��U���N�������)z24^�\X�vB'/W�G/w�L���;�v��2ys��n}�sD�h�r$ TGc�A�y�o�{�ZF~ƴ��>���ˮs�M��Ζ�8y�+��{dUK^���/�&��x�����2��i��u?���-_����*���tm�X~��m	�ȭ'�]�n+��y���,��ǲ�ᯜ�y��@��J���?�P�A7:3�T>O��:��wp�2!P�u��[� �)s\�q0�A�v#C�΅��,-��1O�������ܠ��!|g1�XOz��ժ�W���$�����3����ʘ}���|6��T/��lUD.N���|&��)S<x+���� ��(�^��x����:8u���;�6� ,(Ə�~�x�Ʃ�A�+\�>T�CJvW�v���6�O�c�n8Cy��!��|hr��6���z�D�P��ą/�,��;&�����XZ�[|ͩ�����Q萐��tqf�Id-^p,�J���x��ַ���x�-����}k�s3ۋ�[�_-ic�y�W3�8l`�q7k���������6�:�+3�Bif�?1̟V�:���}���VC>�ZC8�
���Gt�s�6�����d"���?�8]U-�_���jU��ÚB9�x�Gć�����rL���S�G�����D�(!7۽5ǿ��'�Wd���T�]�|�o�=��O��-j%u"e�,O����uD�� Ȋ�o�����[z3)]f²�Ҕ���$x�ģj�i��N�x�za{$���p9ե����� �G��,�X�}�(�V�TO8��;�H�O����L)�{��$��#��¦�t�D����o�#���Ɖ�eQz�|-��`�Y� ����VEl��u$���,��PO���#l�-q�"9�?%W�z�J~�(��	ȱ�����te ��t=��,����9�ږՁ����U��Ӵ�ө��g�t�!���vᐪݬ2
���n���4&
Z~��{���7��Ũ��^�o/���<#���)������s1�����bךP�n�)����L���TO*�_>*v��[��5a^�z�6����������횦��G��[y6 ,i]���Ef�7ϰ�ɛL���C_Voj�?
b��"�����r!��v��Qv�%A���`K7����$�V��(/&lv�(	�˴y�X�H�L�6|Q�k���7���m�M{��8h��Q����i2[R
y�@����pآ��]�I��[r�mRYF�u���<�u����U�� ��-�Y�3��`�� �a��l�j.b�=�#��b���Q͒+�uz����$�%D_�K��0$���� !f�ؖս��B�	�B	2�#���V��˜|�F�9=����Zc�����s�%�����Z��w(�!!�o��[L7�eMr��	������͊�ex��z�{Z"�~2�r(aŽ3��lI�gξJ�����x�J��1ܺ�k"
�ƶ�	�<���	Qև��E�����n�v���;��-"�snS�a���M��PA�SB�^�Y-�u�W ��k�{/@�0������+F��u�y8�C�o��n�J��������j�>I���i�'��� �șBE��U��'[$,5y}�ϒ����`���,B3eq ���U\�9	�,ړ̂%����N�t�N��w7Z\�1Z1���R�m�K72�u�oҨX�J{��1�����7�fx�%��"tX��>z}���)뮍Gͻۧ��nYjӥ�sT֭�*�T v���}쌻��D\5��=�_�_�|<ӡ���1�)sA��ޯ�v?f�ӽ`�c��ۖ�\���`���>~6ױ�j�H��1L�]#y��`�ҥ�Z��sRx^N�bs�������.܏�%o��a$�{��TE�8���jʧKz��"ė��T�,���2٠�����>s�¢
";v�D\NY�e��T��n��j�������Kϵ�XO�(�y^��Tqz��G����#i���pB1�2����A�D|�r��y�� JK�(�n���6E��y~Uz��V���Q�����Pkя��;(�y0`�� ��7������Y��L��B��F��2:�z�V��rDZF� ��$�'���m��u��%pw�a]CU���N,C%���-��ߣE3:�W3�Kq]�珆�?�&�^Fh{{�P��1ŭ6^N��"�6ܤ/{�&�S�h�4xW�(����`��`._�7����a�i�������������e�G����������4�>C��������y��[�U Ѱ�eh���}(eo<�!����朞/�W��q�Cҳ�?�gZo޵���_7R�ݥ��Q/������ᐚ	g�3�E��sc�й�簩ӎ�`�Eu��y�=Ʀ�z�N:�!�|�����Q�ۉ4y��M���x	����ʊ�����,��:e�GE�fi=%\:� Po]��-T��:�ǒ�CKQG����:��.!�����'<S�����eɕ�|�M�x�}�::��	Š��{���1���~�]�j=?VT0���Ī�H��b��YGg;;��b>��Ӝ��r��*��wK�2�;�R]D~�X#G(��וކ3q�lF�)k!)x��@�+Z�\8�K�����m��J����-�=�8�&��q��(��\J�\i��視�������C��x�ؖ=�Qqݒ/\cg] �:��RY�|��o'��;[��«��R�u�RI��y���%0�Hm1�� �L�	A����lS�P$wr4�W��>�~���7w����w��Cgpvb��3��[9�)+.�Piv�U��2�F@W�u�\[�W�Q��~3��bC� L�q<?�,"��U��W�5�>���p�x�ی�����@�@)���\�M]	7�ᵅ��v�=���̽�4�v�0KiH��	c���XQ�{��×���EӉ�ΰ�?d}ަ��ɯ�^���QF�+M�D[�� k���P��*��Hqk@M,1�X�J�E�}Й�����[7�k�sP�<�٦�B��_
=fd�UY|}18%>(����L>9q�v}����e�^�옆)Wo�U��Z�����?��cx��L��u����zo�fL����'C]����=�Iȡ���]Β�PH�4����1O�UR�	�fO�EK�d':��"�O��Ӕ�J5x?6i!* �ӆ~HA)��Q��y�����d{
^߭xr�-i�?D��BލU��7�H�0k�����Hv���c�}���T�g�r����B8v�C#uS���%8od�14��Q�B�'ɨ1��8�%��/�"����u��&'\ �(>?�8��Φ���4�M��@rE�Hn���KL+#�ef��#�<,j�ӶǕ����}��U���x����Kf}]b=��TF���y�V�Κ?�b0I=u�PIc[�J��7��dz�Bԫ&W�ec�.x[%��]CIc��i*6��Kt�v���"Z�P¸بw��yxX���Ɩ��7l�����4�A:'�9T-c#g~V]M��rY@�Z������GC/�߷z�����r����z��"z������O�,�w���WS��M�@�zr��یe.@���Gv��N� `�#$*���;PMv�~�qv����]��b�Ǹ-i����Fo�}�� o$.��������=^�v�e�_~��X!{-��J�v�S�]�ã�Ұ���8Ek!u��9ɟ`:9�0�t6ʸ\Ap�Ǟ0�E���<��r,��	�բAi�S��J�cuO.� D� K���J����|�
@��8SD�s6�|��lMlWN�4S�D�����B/ssRw�ǧ�>��	��BD��2���H���xZ&����1�N $/�.��k�|��V�2�^�Ǚ��$_Ls�j=�!ߺ�_�P����*��Y�Xx�j�F1c4����00H�S�(�����n��Ƒ��1�+�O)ΦD]ʨ=~�O��f�xN?�kR��$
ՊZ�U��5��Xn�'�$T`(U���#K>Ǎ�=J��ށ��<�,��ė����[�x9�'Ӯ�9e��/�e|���<��RdĀS@\f������Pd^�R�n<ʷс�v#���:��r�!ʇw-v�n_q�.n��<q)e�Yw�����;���2B���m>f
��#���ME8��G��<dߜ�n{���]���z����>�I�����*�:���6d�:� }>.<�G]��c`��
�j�q�$h�{��S`��k>W&R!g��r��
	�XU���?�ѐy ��,�w`�҉�������)q/���~�-;���"N�mm�a���6F�����(np��f�cLČ|�ݥ�>��[5���w�X�p�6D��
��z~e`x���C6σ;�Q�FO�hn�N�ɀ�/������W���
�2�V�-����`�~O߁��6��%�Sm�5�g�2��b5����ua7�ܹAR��&d�&+(�(z����3��+<tE��ʚK��b������^|�@��� 	t�ʔ�-~�4)�p�1�TKϟ� �Yѥp/5�9A��CUϬ��P�Ϩ6�%��g�이��{H����T�1��F/��ꝃO�k.'�k$����,{�����.����W0��������0|=�<���,�x��o�+� ����l�E�*��L{E�6�vȕ_`�$?XZ
������a�,������#9�M| .�,i�%�T�Qj��ɦp��2�R�K;_��o�]��0׉>ݨνB�k�I�2�mPQ���m[����_ɵ�<w�A%.|�S.���#  �%J���x��A���)�'
�&�L�r�:�*K�+z�kF��ۛ�Ff`�ߘU����%׿"��\�	�*a�[�.�0��fx*m��_��`��	�,j�167q�����j�(P�h0����S��C�1C�P�3E��R��H��.���6d�w��y���˯Ժ�# ����m�sy�2�XZ�L4��"-{�`eǲm�`v��J�	��
��i����E�/�;�(`K@�e�d'�K���[)QݘbS�"��0k./�(���|�>�N���AQQ�ݵ8l���"�ߟ F��`߁�.W<�e囓�X�ˀTd?j�Y�&�g؅�e����}�_j&�+s�N��j�TH6����Kk�@�\�r�����&�b�������& `�6��
�㉟F��������]¸�S�m��a݄��h�v�If��6�E��	F9�5𹺣w#�ѧs�	��K�>l:�k���d ��pq��σ�i�2Bl����FeD��(7'C�p���t���a�%�!�k���/	��x�� y� 1B!��Z��z3;?CG�֙�"�3:B��F@�Nb��\�9��hd�N*�ӆO�Ǽ.���!�(J3K��{�ߧ���p�#��N�
W��PG퍘�|S�\
��d��ꊦ���<e~�
Z�	��_5�(��3�Ї���=z�LF�����nPQl�Ԭx�f�CnZ\:i{��R�A�]�������}I�E��{�Pu��;�t�ixF|�C��zaH��{�~��JNo|dį2�`4�c0U֏��RA��JmOd1A�?9qiI_xil���2��?F��G�,5��t�����j��/���E�`��L���$9����J]�.�~��E�{�<��$~3�k�F���4���] ����
V���s�b���)�nbj�j��+�7� �6��j]�b?��;�R�|E���A�T���h����䙐� A�[��5����͙p��������������q�R�e��k�+��Kv�Yd�dN���y�ln��N�z��gxj��S��g�D���uv_4ڻ}:
���O�1mKd��S��ͯ�i�P�~�u��"�V[[�M�Ζ��,���	'���� cKc�Ry�����뙋������3�0R������2��O�9t��W8ŤU:�'K�ie��A~�>��p,�Z�Y��a�t��}��� ���<�q;���IW��<军v��z ;1H�\7��KG�W%��d"ؗ���?J�0H5*�0�k��I@C@�֏%C��oM�C1��[:�h[ ƣ���1�0�����Am4'~v��=�M�C�iQ�'���v�g�@����M���B�	���K��W��9.���Z'z�tr�Y�:�oo��߲�����t<�q������
 ���A!���z������@���=����=����W�>��O�YTF�neH�`^+^�:_�D9ܟq�4i�D�,�J�<�&�}=55��W}k�|'�@