XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��uĮ�D�߿��w��2��,j~�T�g�Y��EI��i��1�3N.J�|ô�
�0ީ�]Sݧz�O���F|�5V���9>��ƒf�8@����O�;kS��P������L�^�u(�"����6	��U`]�;�ݛ�ۍCp����� �8TF_�EKQ��h��G_~
���6��M��S���,ȴKz��3dvC�s������L�i_���]Q�68&��"}�w���#�]O[�zz�&���'�m>���t��w[���4mZ� ���.��=3V2g2����<����C��h��[ ^$Z�*��;��43�]� ���aE?���) ��L�6#��)0SU�����@N9��ʴ���\q����yRN�6��D��Q���j��B�"��1p�z��<8�;�i8�U��H���s���|C�a	k���K�JF0�o�o;�S�+k;�VX��ۿƓl�I�^1�i�2��δ0�#ryl�M�oiQ����AI����ss�wrBE_~>I>���j֓Ur�'C������[?2�{�� �i�;�s��+��۠�=����K���<�o��jf�u�=5�g<*�"��j���Z�F���՚��Ӝ������^��+G%�IKb���=����&iNK̃� �7avjg`��M�;�H����NA��NB��%O���/��d7I��H���)b ���I��=������{_�/��|�Lh��ڑJ��o�i����m�7f��~4���
��ßl�XlxVHYEB    6346    1790Ym�[��
�#��s"v>{��X����fp��r������F��B:��;C-4 $��/����mF'�Ѷq]k�X�is��X�
�P����ڻ]F�~D�2ӗE��k[Fb�Z��,@ �O��4D��B�𿈱�sa�8���W���kԅ�P����F��m�c�ߞ�,I�=�Bl�u���5����'	V�$�oz�ߐ%D8j�@L����4눵���GZHm(�@l�����jۙ�qK2X�,�|*�U�$C�cX��&����ͧ����l?qlXj�Ї����|72`{�ؽ]�����Nd�xD�/�7zG]�%e"K-ªC�L}�h=A�vC2<��Tl���a��]5��4��!����S�'W3B i�n�(���.��O���՛�Խ�:�����o���2�w�']��"��_:ǫ-�c�H��`��Yor8t��c�	�gt���~��h?.u�	[�g�4��i���p�%}P���零��:�Ȼj$�ӑ+�u�\P�L�[�HL��<��RP�[��N�A��l��� K;U�&��2ԏ�b��zZ�u3�{v�\ ���t��x�6Kr���m���$;{�4�l�7NΩ4= �I[��z5h�0m�`����q���(��l��J�6K-�<]�ɣ�YфN�[����3ۊ����!e�[�o]Z�*�kW���>�ӏ��]���j�)@�D:@y/QX���{[���g�c��h��\oFckB�J#��H�[z�W V��>BE�1��D��4���T���	���A��o�c[$�����[�vHb�w	���$2���7�E��& �3]����3o�>D����S�
���ۋ����ʸ���=K���8,�:��0�ϧl��^&
�Qr�����dsP�&,z;��	��������~=��&����+��D�v��d6]*hR�?T3 �3�#n	I��e��~s�Tw��|[�����R�ۣ톴'��qT��gmMh���v���ȗ2����0"�Q~�~��:�J���S�J����/�a�Q��?Wnvh�g��XK��}֫A\���߫F�;�<��_��+KJ����з�J�z�%|�΅&��d�\,\��X����i7eD��ѕ�8�F���tp^,�W��tb��ϯ������[����dwU���/M��L�b6���ثiK8M6ޟ1"����؄�\��xL?�C����m�����@�Zm��z͌;��9'8�����G���G�k���f�{^�_ 5ׁ��:el%%4��\��0U̢H:@�f�X51)�l`�K��:�2��d� ��<=�bu\�w�����}�	�*�bΑ��M۔�:|6C�ԓ��tT<�d1[!���%��+;1a$�a}m.т�p�x�i3[/N�r�bW�Eg8����R��������g�(vB�[��=F��]j�Ο[��C|���� 	*�'�ؚ�Ix�v"
���- #���ٶ��Q���W莨7������;�X�{�_k�=#q�v]�� {��!�.��eG�
��!�0��I��FY�	Q��t+56�
<��CL��݆�eӘ���Ƥ=��.ޓ�\$D�H4�(�.�'�;H�``�c���I�HC?���k�����_!k#��g��.y���ˤ*H���9�۽@�[��5u9�V���q'�æe�;�[W�}O�\�R1�1�y��S�l�|c���ү���W�qQj8�L��'叁�&���	�%���u�.�݃��2�T�CH�{��%T`@"�[7v.�p�m�aDr��7� z�[���t��7�@Pz�Dj[� <Z촬	D�8�j�
:I��R|�4@�%��>����۲��x���>��Qm�4��H�f���>�#���H��C�N��k>�p_��")k�#�o���dU�����R���'�_��R0����6d���m9��7ĪNcX�P�?�g��q�~-��������lՈz��K#��Wq���OSG�\�Bx<u�!��.�-{(�(�)Y��������,J&s;�ǌ^�W����p���D<U�(��(޵�,\˪��j�.`Kgj�@.ї4�H��NS p���m�5���=S;@����-h��88j�Z�a���ݣ�1ɺ�G:���k����%Վ\���Z��>�qOP�\R�>���5�R/��y����*�[�iLB�E�*Ӵ� P�bӊ�������R���4Ժ�?���=�o�A\�ڲ�������i&N��ˈ������k��v��Nb���BO�Dw���x7�<C�ߘ��F �"������C5����wdQ�{cN����lVl�Ko/��-6 6ڝ��5�.��f<�j�Yʑ}0�!V�FTJ�Z��]��p��R,��%8~��.�[�������?�3؉jp�N���iP��V@.４���^&���䲕�7e�P����(^�$
׷�t'�wU��ء�]�	�}Aʡ%w�ß	�c�̨�n���%�>z�8���N-}c� ��^۔�Mq�?����7�}13�[$�]�8V�/z)�9��C複dҶ� �;� Ѭ�L�榖�hIE:LY��1�Z������	�$]fv�ĥs՗7V�F�(�}ܿ&��������j?�8h@�~p�Q�u�n
��Zͱ�f��y�H��DOb=����ꓓ<ΊURD�E�1��]�a��*���-�k��a�&D�2#�DfW�I��<���?�0�^jav��{����7��)�9w�}:n��
��Q{]$J��k�(iif�ß-��2X �s�lӖ�b�8}x��^:p Ŀ<yIǊZM�ۇZ��r�K�	�-:��!�g�~O��l��«,R�o�C��H�d�2b�87��be��7�,����!�c.0��0���٭�<�9U�F�?��8����aN��D�rI�"6���;@ e�D����5�x�m�9�'vr��N`�'��T�9#^h��< ���Y�9ɜ[jڠ-����� %.�8N�U��si��b����LjR�<��{��Ƌ���*�� [���ƈul�)�Ob��H���h��q��l�&ݪ]J�y�iDz��� �]ៃx�	(�W�W��
z	�>N�s(*��f�o^<�21PɈF��aM�]��"3"�T����tg<ʯ��U��q�_n<݊�c�D�u��HI��:�Wjm�.���j:���Φ�^\��^WZ������7�a�9�s��ZH�����aUe����w�yO�Na^ղԇQ{h�(�Ȥ}l�̴�VE ��L��2?�.�D�Jes�Gt<��"�'Q1�����ռ�7*�7�K.Dm��8cXuDr���4T#����&��y߫�E�a��{#Zܾ @{Mp��� F���2C� ��Lz"�&ؙ�Kq���c縊�ϵ�<US��!���;��RN�rd�x [���aJ�L���w)���y�u����M�hn)�쪧��O��N�F�(fS���MR9N��*��.��F�\�ت�T5Jw�V����zq�A��,��*��[h�!O �~���e���u|a���B�5�ەrNb!B��h��_с�n�9�� �x�.�X6x{�"?1(Ȟ|2u�{�=J�� ��blw��w�-%�!Wgdb&2&=a���h���`��*;�"�޶F��3����mh���ث�,� h��$k��6P#�a6�!�����N"��O�k��e��ua"�k%"�� ����!��<��Q;EW- ��"uK�e���!���*G�)r���sE��,�a���&���B�A����NZ��5�Z��4:w�j����Hh5��\Y�ILq�����P"I�B ��o��xo�A�{�؜Gck�~���/m����Eȣ:-,n�ň��{�#,>��j۞�fR���T�{���k_�v����ƃ�,+���	"�=D�X��Pne���
��C��pf#���9��S��(kJ5���Z���|�,�!pD��!	�l��yk�j"h��1~�����-�r(������h��6��Q�>��V�����s5����à@�Mv�i+���dU�h��%��S�Յs�PY�+7�iMR�`���i����:�r)����c	㺱p�uT��p��˳m��H�"��j�.�a�A�`1-����:-XQA���4KK(�F@YT��d���4>��������o��n�jLB07�\ g�}c�f6��ؤrE�5B"݌�t����>�q{E��_� qѐk�6�?]X[�&Q ��-��'㶫oȹ̝N�ڧ�+�j�u]�J�	&�����;�R��pL�#����)1=J/�?��f��/�Kys,��9|�xR��T;��z$�����n��f��������t�#)4*���o�f�� RdO��kv����Q:$<���t~5�0/�����ޏ�ԡ�
���?��/�W�}�$8#s��5��3ny�ʹ�EUc�NFm���3ʧ+~���_�%���?���d����j���Z ��M��o�/���P�(��A�/,�;������bUҦ�k���>JtH�P��͘{t����s�
[$2W���B���~�>�P֘7S�Y����!C�J�ﳸ�lF�z�1u�4rM��d�'��m�8r>J�J�Y�׷��+d����}�p�j�#ش ���ۍc�~{kb�i)���q���\��@|� �N&��9[�o�w�E�eJ�A��5��=�PƁ��~v�L��J	REt�����Np1BR}�G�i�j9Šx�,.yA���O���w���������Mu�v4��A�9��x.��\S��0�ާf���vp��J)�x&5��%|`$�V݄v�� ����σ�M�����}`M�l�z���UT]a$��e�i��Rܮ�_uX>W� �����⇭Nf-ZЏ'Iy�*�!��Ha��,��ڔ���b([c���A���+ �6؈G���e��ߚ�۟�����*뮝h�s���	��n(ū�N����Ϊ�r�Pä#���R�Z���HRa�o8���2�B-zݎ�,�W�q<�>e阎���2��)�EFg�7v����=�g�ڋs������uto���t$�p����ֵb��7�{�!J���?+�\�s|�����eV7oIcJ�Ψ�r�(�[�vKG��)n!Y�`c��\f;����F���b*Wǔ�'�Ln`-n� d8Կ��6�i�,w��ŰuC���7�8�5jP�O9��*��FAa�W�žRX���;Y���"�+D��P��p����<*A���Z�g���>AU���G�5�V�*�i 7�~R�-_ňe��R��-�>?i��Ciu����/VN�؄f ��m_����mx�C��n�⛖}25&�HC;K��ai�.�\��1� I �IM��'����)��4eN�v�o\����o{5�	 9/�m���&i�YVkq�Gh�F��&V`�@4�[�$��'ң�#)�L{���nWHZRW���� 3��E����$�dߑ��=����o�c����n2��sWHBupn.���[����;����F���k��'*�+Z�N:��~��KA>�CJuzi��)�m�s�=9��t,�3��"k�s��hO������󦂦R�i[H4���%�����So1zhʹRc�Q�A9�� 0��0�2u�A:
_A-ɍ�=p�a���DH�����z��d7_dR���y����b��`��%~�E�RX�E }��FV��,P����`�n~&PI�E���U@�_�ҷ�������@=D��}b!_E����#�1��H��C�S{}V,47,Ueb�9�U$��Qh����&��)R�3n-CES���B�喨c�VM��jd�w_ˣ3]���Y��+��3�