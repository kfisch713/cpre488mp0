XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$��՗�m�X���fzZK�$
-Wδ��.|
�<�h	Vr�L4�p��_->�W �:��EF0��j�a3c;��_y0@*�Z���ۉ�gsLiB�[�ٮy�w~5���rE�oO}�,��Շ�ⓗ@�}}�:מ.Ma��Õ��skc��W������|a<�p����k�P5�3,.OR
�3%���A5�-�/���/��%ܵ�����V�CAN��E�Ir��fw
_<�[SwwmX-�ㄵ�����g���K@�a7=�ȋP����B�JNP~��x�웆�&�$���/00���x�j�����`���x�AV���9l8�,��k�)k��+:� y�JϬY �D˔3��G{t#�7����u��f�&x=U�&�8g���������Z����Z�<a������
�,�I*��=tdDIʏT{�"Q�A�"�j�0���q-�&��zO�!�@��S��H�ĝZt<d_]"�ﮄ�C�'Ï�a�Z�V���ƀ�SB��I��,��;E��F�N���b�S(��F>׫:���-ZPaFh�m)�b��'\��&����H+�0Wz���]_h2�J,	FקU
�C�3��:ql�]�.��2�o�JNJ:o�¦N�V��0�]��_�Y���łZ����竅�'����įc"X��9�Q�9��\O�b���!'�bKu��5.T�� $W�*��.�$Qإ�;�`]t�yO�D-� �\�o4Vj�߸���)VXlxVHYEB    6346    1790C��\o�H
�+T��܀>C ��-|.z��L�lB��M�jՌ}�>��������Ȏ����?Q��g K��0ϱ����&��]�H��v��-�T"�P3�v�_�H9��)r�uHe�o�_���D�e��cy��j$�D_'��'�o��R�; �J7��H�n�Fׁn%�Ҁĉ�:\l�a�kZhbj���q�=���zX�!�ܠ
�1�ʝ_d�g"�0�IDZ��Z����ef�/�o�7�MѦLd-�g��y#bX��t5��ع8���D���[z�gL53F�@iصR5־�0�D��{`h$^
�W�|%t��$�;�se�C�?�qv����/�@(��8�׭�KOΚ��p�8��|G���k5�f�[�Ņc9��vdj�T��왘*SF��i@���J"�t'��"oͼ��S�����*эW>���җ���*�?�k^4Yd��o
�G��E�CF7u��&L��]:�}�k\8�kƸ4�|�XS|�_�4K�,O�W����m�v)�xFpn�F�"6����4a�`��CyU�F�����$.YHw���B���e0�gl�܁��jRRNY3@��{�~��E���w4db8V-�r��'���P�՚��GC�E����9�'���ѐH^� ޿~�oJ�n�:���F�>t&��C���Z\ZÙl�u������e���"�f�L���>�����1`$�F$��ʊv?��۷��f�f��˭�'�!�׵��85kT5����-����8���"���7H~B`FL�V@�|���#��"e�و�k\���2Q�>�jW;������ԧ�D����͕��k�~�r�E���B(�IS�gQ����0� =���CHm��e��?T[Z�L��w3G2�'�I���8���~T*�?8D>9]�=Wd5�Ъcפ�hb����IF�1���$|�T�����ψ�Wd� $i⾌��C�8+��H $������@���S��Nj:>h21.�k��RV#�v�nӑ��[��7����<URD��p���U���'�X�za[H�S���A��� ʱ���kzئ�H��m��k���駪ٜ�.^?��te�v���Q+��։1�,�+q�5�� ۈG=�`����UCY���8m�����e���^ƉS��m@������3沏�79 L�-|o�?�ń���@B��Ѭb2��&�&�lI��~�Q���u1�G�uT)t�z��8�|���Ԇ����0N�<��~0h@���s!jU?I�� �\Tƣ�ܷLy��ݨ�^)煲Q�9V#�Y� |wNs���ɗ�b:X���\�C+@�\E��j4���M��G�8��⵲A.���G���)NU�3�cSl�|@aO��>i�ߒ-,[A���{e�h����5�����ؗ����f�/d�A��Ӫ��	��]��~���?������/�[�����e� �5P�G�+v�ЍB��P�M��Q���d����g�Kr�|8��`�L��(��oPe��'ج�H��1�B���J:�w��:]�O�{و��n�b�!>S �h����Ɋ��1R�Ӏ��-L��T
��`���d4/}"X�nR��6h��V��s��A׮6����M�n�����<� �	jIE��D�&M�c-t
-� '�뷾�*wP��s�/���#�XV�D��#�d��p��}b-_%D�������:L���nE�GYv-��9�CNB�	��~�3��ȕ��@8���IЁg��H��oirKdy���l�?\�c;Ǝ��� j>)5K��ƳP�hł��� ��`4������V�nf�J�~�c�qt��,���0Γ�d��@a�2����޿]��_u�����>�Փ�����Z��2:���X �z��1φ���a+K��H���-?����C5�Ř���z�F8�����Iu��;�͔���j����3�&��6,�gD�1�+��>�4!��t�ܥ����-��k�;�+O��ж�Қ�2���ث*�I��.Jk��.n���}������)_��bݠ�0�EdL�}
4~���B_?+w� H}�sU�����2����8�a,�R��v�yQ0��b#2��\	G?}^�$��f+xD&�*���j�u�0�X�}��Vz�Zwup�
�=�8�������I�F�U�kՒ�f�j�pKj:# ���f�|��2v�0	����ѯ+�4:Yp����"��\xVh>33B�(cqd�y�bC�	XV#D�ER�_���2H�df�D�Ũ�g��%�Q��Ʀ ����Dv��d%p����Z|c;-�I&
�ņr�i�LAQ���K�#}�+]:$�ʧ�+��nM�j��T���L���Jz���'�>�{��F����^���Fᑲ�;��]ʌr�u�÷n�����A�!811K��+z���S�2���ڳ<nʯ�����4;��7$	�{Id="�$34��LC�0F����e���y1S���]�e�o��H�p�����.	t��5��HI�]EK�!�A�.�Z�pq�2����"�xH���!��AY�/�� �
���&� ��4�,1����S���c�1���U��?(B77$v�"Gb!I��}�I+��_�OM����u����y&4��"F)�L��_w`�~o!:>TӏN�)7�";hi8O�Ԙ
qn�4�wR���U\A�[�'�iǏ��pj�� WѺ�1�"I�!�;��!�].�Jt�i_�vl::X2m���o��`0��B�똪!Q.�h�T;����)��n�Kxs���I.�pJ������+?���ˡ	�[ﵐ����q��p����%U��ߌcE�%�vh�2�~�[=��t��<&� �4f���a�R7gf@O\l���Q���S¡��GJv�mx��I��F!Տ����2
�̓��"�Ka�'���v�銾�Y1u�ι��`?�2��& ){n����~a��C��[��:�7:.j51����ү	s}���a�K4�kӏ�S�p)#��3��m����M�d����������D2��R�B���~-����7&���k�?*�ߜa�̎�j�e�[��}tn��ʪ���d��`����\JY���9�
���\��<l( ����o�2O0��Naz�����zp���pM�����m�#V��g
��\Y��`��ϫ)|�L���Ā��F��K�
�3Z4*����.�̻���	v=]�J_>�`��8Z��|������/] ���B �)�����9�g;��e�^ /-)�Xۤ���w���QBJY�JG5�㱴xޟP	Yd�I�p���m���Jg�k��-�ޟiG�jW��'�����	���.Gpc��\E�55�BL���-������&�p�Q�7����G�y�N�a�eaC��~5�}����/�ɍt[��V�[�O�}���)�ut:+��� $w:S�l������,J)�V^�M�Ƹ�<�� k=m��>}��]!W˴�+勧�vv������"�����įA�S2�������8���y��E��:\:��R
\�K���s��nM�Јw�G��%_�ow�s�L�S��}Em��S�G��o+2R��h��X:^oFyp��H��2�,���)�?��Z<��f���}Mf���� �Ʈ�oI�����Ɨ��G�v�՝�e�v=���1gZ,c<��7�j7|%��l0Z�*��nC(
�����)��0y8�m�����C�`�ś7[�'7}Z##V!��(�gz.i�����cH��u~a����Ff��i$�	�N�v"O
!��$�~R�č�́}��`�y��x������4�4��>h�^l��!7�d�z�$:o�(v?�����d(�&a�鮉�H��r>5�o���m�����x}�a��-O-i'b6��*���s�<#�'XR{<͌N��S��h�ul�a�ї�b�x�2�j�֓��������!Z���G�?|��yq���rzG�JZ5��qk�8���6OL�����p��<�ت���r�N�ju��K��ۂ�OM�� ��7�����O*]�Y7��i*_�.��^�'\���!�Έ�.���f����VF�V ��!a�G�sd�).),Lq�����ʩ��?��J`SD2}�g�ޥ��`d��r`���4�y j��>N�]K5e���t�e0`H�#݃�;�*6F���%=u��r�{��x{��I_'�m>
v,��9݃4�A{ �~��V1M%᭫Tʳ�u��b"�Z3R>U��,:����<�C4�,��b�5��_�E)n�v��c�.��+}χ�$��(0��/�i/o1�s�jL@����'_ �QZ�7D�b\�|�m�_��&&��ڕu(g�*�^w*�M�:P��)��ѓ��t���ȒN��sʅ/x_o�B�a$C�gx��B��m�O�ͼ,:�e�G�#��B��b
��ב������H�nb� I�#�h�C}��޽%U���W��WyEf}�x��X6X�'�-�+�C�3� �L�`w}��i�f��L�nC_��j>u��P͋AeR��sC���GGr�;ڎ�&��ꧨҐ�rW����g.�).���i��|�*����Cn���_00c�ً۬1�;L�����"6`���4<���� ����I\��+����mz�8�Nt~Q�F�wB�������h�ܵ�з.� I�R��Ur�
6�ȒM��h�qd�P_a`�&U4eV�15���&���V��F�l詏�%��vې�^clSgi$6�w�*��G=��U�b��M�]�4J�nA}+�����3��i�����PE��r(W�"��㪤l�R0�;D4��5��nKOpX�3,T�2P�G����u��v����"��m��ڵ$��&���Sʵ�v*ć=��Hv��fO R��U��Nt�:�j
D��c�po�;"ȟ��р B��\�Ƀ�`�,{EWOq�w�0��������|��Je��U��`ڌ�P$�vs��Z����M���|W9HN��V���;,)+l��Q�ƶ�{��׵�7�wR��Qh�V��p���U�m�!�YC�zi�RwN��H�q�}���+�|J?�f����=�{�!��с���oӪ��h~�u��8P���UG�M���%��Ud�ߑj_��l���>Da,��;#�H��'�x۫���GUQu���X�k�B���2��r\��4���}���,�S���/�By7t4)9n��Fa��b���tt��o��>@��:|ʸk���N�'�=��5��R1���4��XZ�6́)I���� �����]������>����.��-�uj�nW�P���M���D�9-qR����G�rKH�jA<��N'I�@��Ɨ�����d
G�� ^��E�q0S�d�3n%ƹB�Ә _ș!���_���D���n*E��;��q���i6��c��o*�n���oj	Hvm�xe@W"�%��;�@#�)��Ծ�Xx��e�k/8�H�o��Θ�U�T�"�T���#%�5'K�x՘OW�
ф�z�@a\�Ӯ���(G)|f9y�7�B�������I�~ �!�8� v�>��PK�h	37����)��G~Q�k!�ϸf��0��[߾HS�����p�w�V��̬%�K>������qu�+�r��ϥ��)��&�ޮSt�'��侀�&��r)���+�3����h�Z|b�I�'�]:��(�!��u�E�(���w$vl��o\f�@m�J0�<}D[��6��e�U��
il7`���ڽ����c��9g)��j{&��z�x��qc�.�o����o�N�+�bb�����:�Ѝ]t�*цM!�����a�[f#s�6�0>
<��%{9xi}`ۯ��