XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i�?��{�I[SvW������uN�<w��g��aC�w3��+�nn��{�}�8FU�Po�M�4��3�8�:�������eu:�h<�2�ޢMr��3Ԣ�6��7��~�{��aB7�tO=ϒ�f�@�#+eE��T��s?}�۽|���`|]T�;v���ǌk1ݓQc>��ˉ=O���YMduh�=����O�]���[P�����v�t(w�T�+e5�`��9�8#����cDz�%�N�k�n����G�žÖI��f�I�Ϣ�g�����=u� �I��g|���G��5q*�]�x�XT43�w_�w�~�vm3���f�x
�GD�ڮ���bU} ���7]�<13|�T:��\Q饤�����Qz��5�����S@+bCb:ܚ�����*185h�j�A�s��6f~��d�ɧ�~��`�wƋ�'���Z"��w@�3͈V����O�����UO�=ń��Af��;X3P>oD�-f���ğ�j��H���Lz��vٰ�(s��͏eϫ��<�{N�7%��#�S!��̃�AOp$�?�|��OB��R��O+�l��6|�Y��o�)�ޤ1W��B!�YhQ�ܲ�W�W��.5�Ӻ�����M=�lԲ(�����R�1�D��e:�3Y� ��=>�W]x^ �{6��ӊ�r�{9���o����b���C|/�Q��V$F�T�j� 0E���U�	ϱ�?g�5K%C�����%�>)l����[A�$�������XlxVHYEB    6014    1840�8z!�/��zA��,:����8|� ���!'�,��!;[�4���)�%c6^��,=V�2�# �[[n�ą�gt��b�N����J�GҒ��Yb���	�@ؾP!]�4j	�˺�P��()�3\|��aXi\�͈09�D��~�F�	���
������4�5��
��R�� *m5B�C�^����?߲r���X���Z�\��c�{E�.�R(�͏���0���&�޳C�ƝF�"8�#����}:�����CǄ�odl沦�5�S7�`��7�W4mf��~���|&x_0��/4�Q"K�c��ͯFa�/�L���@��q~���H߶�B&K�%؏����UV_��y(O�Y(uߕ��"3�R��T{-gS�R�X�X�ס"�HsoM{5�vuTs}���5�!�y�c���O�Jr�z+��,6�gh�ّ{�"���(Z�3J\�����2�B� ����Mi@.�3�YaJ�� ��N��v�(���l8�{�F��,I�8	/"y��y�Jp��G�o�%�6�Jd�z�'�kJ.l�F`��T�j7����o�+-��}��zE�(��A�I���T<ԧ��e�
��O�8��6��B�������J��pVҎ�<��q ��O¬�;M�=S�PȾ�/��S��y�4���	��t��u����b�7�w�Y�xM�po��DY�۵C����i�a�M�	s�o-���MBh��_�A��x�����?����׿c�+��V�H�PڸC��be:xF9\YO��7 ��So�I2�$:h�IW���C ���g���-��l9(e�&(��PKnyX�s6����Oٰ=�o�hnns�`�}�ꀰb��l;��.I���t�L&��c�Tx�Y��I��I��\BK!9T�(;בs5�M�S��x�ˮ�)�fM�h����������NRK�`>f�bq���]��;Tpfݨ�K�}+RE4�!��Y���@��&�.�e�'J�/H�Y�������$�ݵϺ��	puW{���V��lgD  U
=�S��T	ϛ�_q����D��QO�㿜�djD4JC��;�tX��(|�x,�N�(����WL:�xF͟��,Zn�&k	���paa�y�^�u�'��'���c�+�G-'V�8�.�n&2��qY�Ψ�v\F���&��z�c�ڮX{�WjO=�/4����	������7��1�Jv�X���[j�>Ouy�&[�Y��gj���H!6����WZ2���0�\b��{�T�@�8����Z1�<�:��䨵�~◌�pu�y���Va���Ϩ��bNgW�F[tl}q/?��s�^��������^��� 	��_8�m^�r�@�-B7`��� �G~��8���9�c�����T�ڠX>�;8jE�@���lYF4fI�9�i~j�=·�H-ay�G��a�Cu����Y;p��+%�HVT�����#��Y��$�F��+)�Q��F���W�����eX���~�L!㴇@�3�FX/*���O�^��{�2�l�6��&���%<(_hDˋ���)�ڨ5�����^���x� ���`��V�UD�n�M,��>����Dp��\���G�{5DS����6���he9d+!��Kۤ[�!����]����;g0R���p�n�DA��Je�&&ǹ�(	�7^�ms���4��/���}@а[�ܟ+��D�դ�gu��E�^>hΟ�30�`��RB_Шwؠ�OT�Z��A�go#("�.�_��w8���5�OR���Mx�P�l4Aw��%���)�Qfv�������S�E%�"_����!����r��h�QX����֓��6�t-^�5BT�᳥! *��\�Ɛh���G���f��dq��� rJ��^^��l���*���h�[�E&,NwZHC��p}I�i �3}.�M��=ƽu�ߐ(���c����K"[�}���z�T���侟��ݞQ������|�3�7��#���(P�6��r�����Ja�	�8V�[�bN&�����	�h�4�JP�,﹙��o������H]��{2E���QO���gq��6I���;&�b������7Y0B0��i���o�u!%Z����E=[�r��N���NB>��nP+W&�Ds��I��8�J1���V�Kn�����gΐ�n�z�Ty�d?x*&\�ʠk3�=RR��Q��?,4�	���%W?���d�~�\`�:��xv�v��L���<8�>|[{�`4YYb5���m�@}�����Y�{��l=�=�BZ��~�X����h�ڽ����z���Ů�N�" J�����X����Iz������+UT�މ$M��ac!���C���U"B���q�[[�e��U�y�^MWL敍�v1���� x}PiM�x�^��<�"1̶x��'weV"r�LK읡�cJ��K�hS��d��[����8N��d����5%l1\���CI�l�q�m��
ߔ�x�L��|�m{�u@w"�_�m��W<�mti�ߜ9o��`�n�J;�s[����c?��)�uc.�ećm�u��a鑯`@|2���b����Mn��c{�շ���JAyZZ���K�#�c��$1��9�T�BSz�L*f�m3LqmB3��A03؋}G�L6�<�z剚M] K�ҷ3t�7H�eD���V
r"I�7{�E�m�к�p��W���S�Ŭ=����R�<|��\�Rra��C4KD�����)�炩��\h��sM�Y���5�ԩx|6�i�I�vv�'Ds���3�a���o�A�1=��|�Ս��7������y|��8�7W�Zh�o+>�A1�c�X�x��`^�E�^��c���Ý�����yJ��0U����"�^O�=�a��Y�a����-ؐl ��1O:
+.���ژi���x���3Y��N��wHQ<51p�A�$&}t1-�qɗ`�Վ��`�hw��_}�EI_}{)O���Z�Q۱���P�A�o2���x���n+/9/�zRJ����x�H�E� 4w�%!�I��N>;u��p ���8=b=��3���0ߓ�0Q�Ȩ-�?�v�쓃*�����\�� ���L�����ٸ�5���$�.�ތ�3y�H� �<g<�:*b���$��z�fc���~�?��m�RŤ+�8d����K���n��<>B�������N��]]�F�9�t!C:�ۿ�F@s|��8���U�P�R$�ݑ�q�x�9�.�Cm�<�Os���Y�P��#�M��|�Oo�h$�[��`q�?�&K<�\��g� ��O�b$�z]�Y
w��ɬQ���o~�{��X$D�?�m[�a��fk��yJO��lb�i���ÖN�N n�6w"��ۿI�Z�0v0�yn����o�"���'��.\�Q���=��-G�-�ld��;�)d��O�.t��d4#�� i<yM~�]�h�L�$��l�C�l�4�%��������0���B���@�UX=�`u���A���yul��}�]��(82����gǯѓH�ȒL��$ӤƊ�	F/��AM-�M(b�֢�3'�2棌����1M�h��4��S�2�_��)<)2�/tP����"z��޹גּQp?��7�-��5A6����V��.���*��י�1b���������#��$r�����7�\�ѩ�ȦI�I��`}��H���ƀ�B� �^�6��p���r�?wB�b)H�b�P�G�m��[p���#�"�3C[~���P#CR;����"�54gɐE
���,&��W��~��=��ߪ���6 ��l�?Of �iFo��֘��ߎ_K�+6 �l�^.��!����^iw7x���P����^��ǡjK���OcFP�.����o]�%�j5bCJ� �_�t�B[T�0��dmY=����C�Ա*qW����Ju��on�i������\g�}���UK�\�a� !�� ;��~s`n#�Wh�!�Dz�:V7y��=���?��!�-����Y���}��s�F�r^��mՖ � �W�3B�������O
�����]n $�ں�t�	��SҞ�V��o��D�<������^�[�.�^�O/� &�p�q/��Xi�e��߯�1]}���y�|["���b��?��7
j�W#����a��މ!x<.�!0X����{9���SQ�=*�3�x8&G��~i��]�$��W�	?Л����nH��h}O�s�����C!�0�Z��-��Y��Jmh�ߔ��(S%:��L��i�	��1P����7\d�d,wkP�B���.�Ɵ2Dc��}�uP��2S�1�q�Ťh�7&i`i�GIy�e�16~�~[����!C4	q��
����Z��ѡ9;������^�ɵ]�~KR� ��X�ʍ4�Cj�+�'gH= ���Q�Ớ Υ�0��VS�� �zSJnm�a	����gm���:P+5Q�(�R���)� �C�����6w�Z�dю���ȕz��&���3T�9�ӝ�k�8��Ž3E�+wh��$yJ����Z�]���H�d�+%.p.��4#}g�t}Wj?氯+L���,�>`T�����T@�����fnӛ���S~C+4�-)��`�����������sYZᩇH�M�<��ɶ�8�(��ǯ�x�Ǯ!�}T�����E��sɔ�d--\{�d����{�bn��E_�h<k����v�:5�[p�����Q��ɜ׸-*ڠ��#h��m��ں�U�B��xƅ��������G�Dg�)Lm蜏ķA���]�lZ^�(�`��g#=�X݄�-�.ռ�&�QO�7/�OɈ8	m� ��Z��h]+oA wˊnyeA����ْ�� >|�m���n�L�65HmO}�_4�T��Cϥ�Kl�8e`s�:���A;r&�L�� l��L��՜��Y0�vs����[07��/��x�{8����Y�w:�ˤ*��P��?�kQ��|���2g�:'����ӄ'��3�ª�0�3Gy���mȊ�t��}��_�F�7�I��J�v&E�'�?H�h��l���~|@���d�V��g=a�x�h���h�Nq+߬�煰8*ũ�5�E�'�j��J��2��Q�t��k�Ě2���Q���J΃����Eޙ�s�Ӫŭ�������F٣��"G�E����h��G_�T�،,���5�u-X����&��_Tw� W�O?���>�՘��cN���.�0��s�b�,wԏ-��"��Jm��3�R�W�&��b*�zvH!&��MR{��#aTƼ�,������bc�V}9��K=�}���Vny�%�<bW+V}��C� "�I��PY[�m���e\�H�P��+��3~��K��^G$e�X��SL�Vr���2'~k��!V�]��)z1oW�9��#k������� ��n@ۘ7�r�T\a��G�������#wF��{q8�
I�� d��Za6�_��.��s���/�����U�|Yw��&a�@�d�MK�U�����Z��I@n4^�l��9�E���(v$��_��j%�p�%���6�#�h�}��d#�׵�ߛp 8���5���(z1ob�CL�m�m� ��"�����������Xd'����D��E D�0Xm�M�^��U4�U�����J�>��X��j�|k�k�.�@�S�-%}Pl�c`C?�O�[",�0�ך�oU4���W��ic��in_5�1����Lث��2�w�u(C:���%�Q+"�[��?&ߧ�"	$Yj2��Y�����m����%�,S�K.��K|�2n��~� K�+z�(�j����U����D
�Nv���6��$�F]c�Fޒ|��י<#��:�����Lz�������wS�]A�y��Б;�����:�K+*�5�]l@GAF�)��!��CZ�bT��Z
.95J�����4����R����.��(��fX�o�xBe��]ϘUbd|w���w�#�,0&��.����1�_� ��"'�(����'��v��c�{O��/ۅ�Vj}C����js,no���g%+jLW��@�[�