XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$�^:x��1��t�O�_H����`0)d{@C�Y(k��:��oYq��������A��'M�;D #�_m�|������X{:�RQ�証����v$�x9��ļ-V��Q��K������1�E�aȷ��+H�����0��蚒�1do��iwף�Q�jڢbnd�3�:��pؘ]���鰳v��B��YǓ2A��ַ�g��RB)$��v{Ω_G�{�����Edk�X�~5�:4}����F�+ �U�+��?����*	��?�Q�ȇ�!QPag�{��D�{�<D[����Ey���7Y�Z9U�~���g0by����6؎c�p�{�e��J�Ji� 
��C�w7��E���S|��b�;b+9�ɔ����} Dwpq�Jځ=���@���7Ƕ5�!y��3V�=U�YO�G�1�r��Gq���	�0�?�E��;Z㿰;"%t{���h�f\� �ґ�tZ�-�7,8J�ė�}�/�EQGx�Y|��a�E����6AU���}��nI����G3-ڨv
�0k����h{�
/�+�4��6%f(�7�1��R���zx< Keڝ��{�@S%�]�_X�(I]
�\�h��x����;{��>�׈�pbP�|t�K���ȅp5�m[C� �PԢ�J��:�h�|?]��c�*{ ���t��AHB���;ʔV�ߔ�Z��(>+0s&ֱ������J`OMZ�^�hQ^�w6��j1,;8Zs;EXlxVHYEB    3fdc    1160� & �b�C�(:�'��$(��'.{��AX�N0�d
�'/9y�P� !Þ�0*H����1��ټ]I�WřDBӠ����7Q�&ao ��vx�V ��х�M��0�8��R^��n\���+�ȕSEw��EdR��q;�-P:O�O�)')����o1)���ν9a����<^���6�t�^/:� �p�%YLIc���7"��21��ލ��Pü~V:���R�vW���<I�┅��(�ɘ�ውE��/�'HO�,��-� �	�N���)�!�t��&ޫ�o����xWG�
�-o�n?1�<��X�6����흉x���+������g���;]/J:]��J�"����ʹ�ժ�V��mm�^y�����I�ƈ�)�J�S$�y���z%����R�Z&,�0���qt����`�l����+F�L�<v�]��'�n�,�7���%IV�Ǒ�|[��A�߯}.���������
��R��Yub�s��iZG14��w��V"]e���K�%��M0�f�LGiEP�wUCu)9p�b��gc��o�Td:��������SC�� �w�����âm�?�Q_�:�7��m��n"<5F<z��h�C��^�7?�W�ƥ��J�֋�G�O$Y��L4��p�I�{kr���u��Ԇ�bU?!~��[�+acl<��А��~ث����aamX��Υ@�m��㱴:�9i �9=!�O��V���JÞ����>���%@���/FV�QrV��UHU�a��w� Ѐ p���?���C2��e����'b(����#�1�Rӆ�.T��y�4�Z�`S�?޽<� ��v������c���k��<6�<���-�瘏(֯yX�r�w��1����n˟�������xOCm<j?��0r��Ԍ-Ƙ!��CA/��-b�_��� T�Coa������N����;AB��jP��FǤ�>����j�5������0P��Z�{��v�8�(�C����l%D�?Rʛ���6^gl�헴�~+/���ʸ2��6\���,Q�p��:r�0}����b	�R�p�4)8{�>�@PM���R� �����E�O�� +��^-W�dwC0w��B�c.w��¡u��Up�j�Il2�s^���"�	�6�+��&k�f����3z�4��ݍI,���w?}헚��Q�:�7p�L�����#u�z��d\~��i�')�y!�`�������M�D�Ƴ�+ �k�����<��AHWI��Yz�=���Px�A�] ���[���{�\l/WI�XN��'q�:�d�ߎ�-`�(W���2غ�ʜk{�q�љ������U�ۮ�"�rz�_z�"�sy���*W�f��J�����M�s��|�U`#b��e�����'�L�a��l��j��3ZLl��m$����w����� *yIc"K�W	��BK�|e�x+^�a�f��/�.։�>v�o)1T��*`&�G{�|�< E:�����H��� �a)�<�pǉ��4d�����\~������H�m�(��T<�R�c�T��M�;Rηz�\'2������å�&=�C9vJ�H��H�D�9��A���5F�!b�Dq7�..?)c:���!N�4O�d���?��R��V�_k7�����z�:����K4'���Y��AԟBhL"��
<�B���0��z!|�Q���ӓb�|������|Sp��O2hP�E�6�h
H3��ʸ+��Kxl�& DGѽ�Y?�37�X����3�i�S��b�ѕ�zJek��oE�q�Y�����iN�i�]$1�T���fO���ؗ�e��˜,�q�Ԝ�C�3�����ˎ��T��Gka ��H��ڥ6 zי7�k�	���9�6���eR�'u��u�o<��m�:�-Ġzz�K���ނ1���nNu�"(�o���S��SRS���E�A����\D-��t�� D�`��~�|���|��Q���-`���t�K����u����
�+r�F2��̯Z�M�7��Q���Ӊ�;2���]T��� ʦ��m&��o	�}���i�Z�'	D��X�Mi��\P,76˳`IU=�(��l�K;�R�����;+���V������!H���#�}9��n=�������	k�3HY_4�vw�!���K�]h�D�×���'<� ZY�KΆe�1X��Fܧ���z��� wLZm���*V�Ԣx$���o��l�ˋEf7)�cȗ��RV��-���̽?pF��=CH�!�H�@+�����7���Bx��Pb�R�[�1\Ξ�ZZd�l��N��gį]VyD�o��q�.� ��sЄ.B����|pN?�2�RޓQ�/��l��N���?l�(_?�_ύ��(��DV�%�O@K#�	��6��^n�h`��i�e٢,3��A��ݾ�9�)�\hڀ t��){��t>���{4L\@�a�լ�b..���L�t8�Ũ�t�.�c�<]��V��.�h�����%�)�i֊f�\��^L�u��8h4���.���k�I�?��@;��#��.LnJ(�đ��o���"���]�=Bs�A��׹`��m�F�f#�������l/�,��T"�5j��(��>����CͬM}�`cK�S�x+nlc�o��57�`��hl���r��:�ȉg���nXɡ�5㩬1�[�T�J����4Z��=��$o�mn1��,�/�P��-St����t�1)����9�KARd @��fw|6d�_�8���u:"sϋ�~�9^�7��#��mR<��d���'�~L,�w�Z�ma�)}��9;7Y������=6x5�cIGrohz�C��  ��CiK��Y��Ȧ���!,�Z�U�.��%�4��{rs7B�R��rT[{��)j��n�i҇R �M����	u^dz�	h�g���W�B6���C��V.����s�I�^9�|!	�a�a`�_-����#�����`��x�q*B�Ļ�σpO@}�C���q$��2l;Y��E��f�5%��ζ���zdcXݓ
���(� 󥳸�(flVg��N��+~G���a��L}���5��"|�����!����s��6'�W�{4�����v$Н\=m�k��.����v:�>��<��7�cl�E�T�k�iV����+�A�M��ƣ�~~����r���Y5"WC��β�P�VD�־��M�l���1g�z@	�(}����-_-��ǝdzp��u�SX@u׫8�h�Y�0l��td�g�3u�ML���{aIp��ES	���-�G��x�T+!��y�Р��hv3g}jk0�_�v��$�d�$��H���8�臇V1���6�['rC^J����]?�����(Y�t��ty@%�;�Ql��Q7��6*�� W�&
���d(�>�gc#��D���h�q1��c��SpN�{�B�/Գ�j��J���٠�L4�����o�X>0��	�S�/^�7�����nȱ�$t��nR��|��&�l0�V�3���q+ĩ&�\Z��^2���W9^lo�����6�F�(F�#���v��_�h'�������8K'��I$ �W0�-fm��Pp���6?jxRku�������]���2k:�j_�ӛ#���I�ԘX�}6ϯ��I��j>�v��v���u��w��آ{���\Sc@C�RMO6�:�����t4{�(e��ʚv�3����X���é^E�bt{+��C�-�� ���2v����:X%�;N��>���;��@I���y�P����
(���uq�M�������.)|#2{ۑ�A,ך&�%~X[r*���i.�36|��,3�1�(~x�r>���,ZI���+��Y{6�6� �|y�(S�N⡾A=n��Qh��W�V�9�Ɵݨ�By����� �W��a��	ʈVK�6u���"{��=N��P�74�Ԇ2�=Ж��&RR�]���q����,�Yu��Y�ʙI17k��my��
���t�=V�bȯ��(-zz.��A��o����<�p��W�"5l�m-�2�xU��v8\T��=¨d�>,� �N���DQz�~"���M:F�1<���tn�{���q��ORj�Xbߵ]������6�b�P'��������~|l�2��8C��ֳ�uܚ�P��T	�,섕Z��7�|�Z1�q��́���W�G6�z�W�^W��>|%둱q��,l}O�@`��fjK4��=�5`�/�vz�@�c�_���G����zz�FD/p�eb��^�L�Lնsks�i�F,(o�YL�X��md� &�V�����b�_�Dz��$X.M�ew��T����4#Ϯ�I{��B`��